module rect1_rom(
	input clk,
	input [11:0] addr,
	output[19:0] out
);
	reg[19:0] q;

	always @(posedge clk)
	begin
		case(addr)
			12'd1   : q <= 20'h19dc4;
			12'd2   : q <= 20'h08a44;
			12'd3   : q <= 20'h09de9;
			12'd4   : q <= 20'h29846;
			12'd5   : q <= 20'h394c3;
			12'd6   : q <= 20'h20189;
			12'd7   : q <= 20'h32548;
			12'd8   : q <= 20'h199c8;
			12'd9   : q <= 20'h704ca;
			12'd10  : q <= 20'h3a0ac;
			12'd11  : q <= 20'h08643;
			12'd12  : q <= 20'h0a222;
			12'd13  : q <= 20'h81882;
			12'd14  : q <= 20'h2c442;
			12'd15  : q <= 20'h708cc;
			12'd16  : q <= 20'h2008c;
			12'd17  : q <= 20'h12e48;
			12'd18  : q <= 20'h29d42;
			12'd19  : q <= 20'h7aca3;
			12'd20  : q <= 20'h28d49;
			12'd21  : q <= 20'h4904e;
			12'd22  : q <= 20'h1948c;
			12'd23  : q <= 20'h21585;
			12'd24  : q <= 20'h29948;
			12'd25  : q <= 20'h400c9;
			12'd26  : q <= 20'h4b028;
			12'd27  : q <= 20'h01e86;
			12'd28  : q <= 20'h380d1;
			12'd29  : q <= 20'h480c4;
			12'd30  : q <= 20'h284c4;
			12'd31  : q <= 20'h604d0;
			12'd32  : q <= 20'h01648;
			12'd33  : q <= 20'h43d44;
			12'd34  : q <= 20'h18488;
			12'd35  : q <= 20'h199ca;
			12'd36  : q <= 20'h104d0;
			12'd37  : q <= 20'h04a82;
			12'd38  : q <= 20'h43483;
			12'd39  : q <= 20'h4b843;
			12'd40  : q <= 20'h03126;
			12'd41  : q <= 20'h29c64;
			12'd42  : q <= 20'h48c50;
			12'd43  : q <= 20'h199a8;
			12'd44  : q <= 20'h60d02;
			12'd45  : q <= 20'h4208c;
			12'd46  : q <= 20'h58d06;
			12'd47  : q <= 20'h384d3;
			12'd48  : q <= 20'h480c4;
			12'd49  : q <= 20'h18523;
			12'd50  : q <= 20'h43d44;
			12'd51  : q <= 20'h00cca;
			12'd52  : q <= 20'h191ef;
			12'd53  : q <= 20'h31506;
			12'd54  : q <= 20'h2118a;
			12'd55  : q <= 20'h31084;
			12'd56  : q <= 20'h7ac22;
			12'd57  : q <= 20'h1ac42;
			12'd58  : q <= 20'h82c23;
			12'd59  : q <= 20'h1bcc4;
			12'd60  : q <= 20'h31d02;
			12'd61  : q <= 20'h1ac23;
			12'd62  : q <= 20'h30182;
			12'd63  : q <= 20'h4b843;
			12'd64  : q <= 20'h3bcc2;
			12'd65  : q <= 20'h01486;
			12'd66  : q <= 20'h23182;
			12'd67  : q <= 20'h30c29;
			12'd68  : q <= 20'h54462;
			12'd69  : q <= 20'h4a442;
			12'd70  : q <= 20'h398c4;
			12'd71  : q <= 20'h3c462;
			12'd72  : q <= 20'h54463;
			12'd73  : q <= 20'h43062;
			12'd74  : q <= 20'h48cc2;
			12'd75  : q <= 20'h1adc4;
			12'd76  : q <= 20'h0aa44;
			12'd77  : q <= 20'h02863;
			12'd78  : q <= 20'h484c6;
			12'd79  : q <= 20'h41c66;
			12'd80  : q <= 20'h08249;
			12'd81  : q <= 20'h62846;
			12'd82  : q <= 20'h01668;
			12'd83  : q <= 20'h380c9;
			12'd84  : q <= 20'h28cc1;
			12'd85  : q <= 20'h58cc1;
			12'd86  : q <= 20'h2a886;
			12'd87  : q <= 20'h58cc1;
			12'd88  : q <= 20'h21186;
			12'd89  : q <= 20'h7b046;
			12'd90  : q <= 20'h48c42;
			12'd91  : q <= 20'h48c61;
			12'd92  : q <= 20'h0848e;
			12'd93  : q <= 20'h48084;
			12'd94  : q <= 20'h3942e;
			12'd95  : q <= 20'h98024;
			12'd96  : q <= 20'h294c4;
			12'd97  : q <= 20'h4c862;
			12'd98  : q <= 20'h44862;
			12'd99  : q <= 20'h21586;
			12'd100 : q <= 20'h1b046; 
			12'd101 : q <= 20'h5204c; 
			12'd102 : q <= 20'h3c862; 
			12'd103 : q <= 20'h480c2; 
			12'd104 : q <= 20'h2ad23; 
			12'd105 : q <= 20'h480c2; 
			12'd106 : q <= 20'h08645; 
			12'd107 : q <= 20'h40084; 
			12'd108 : q <= 20'h1b023; 
			12'd109 : q <= 20'h438a3; 
			12'd110 : q <= 20'h2914c; 
			12'd111 : q <= 20'h4992c; 
			12'd112 : q <= 20'h1098e; 
			12'd113 : q <= 20'h21d82; 
			12'd114 : q <= 20'h390c4; 
			12'd115 : q <= 20'h21568; 
			12'd116 : q <= 20'h1aa04; 
			12'd117 : q <= 20'h00202; 
			12'd118 : q <= 20'h394c2; 
			12'd119 : q <= 20'h188ca; 
			12'd120 : q <= 20'h5150f; 
			12'd121 : q <= 20'h1b906; 
			12'd122 : q <= 20'h70842; 
			12'd123 : q <= 20'h0a8e6; 
			12'd124 : q <= 20'h79083; 
			12'd125 : q <= 20'h125c6; 
			12'd126 : q <= 20'h29d44; 
			12'd127 : q <= 20'h32508; 
			12'd128 : q <= 20'h70462; 
			12'd129 : q <= 20'h09082; 
			12'd130 : q <= 20'h5a848; 
			12'd131 : q <= 20'h000a3; 
			12'd132 : q <= 20'h11648; 
			12'd133 : q <= 20'h31826; 
			12'd134 : q <= 20'h98423; 
			12'd135 : q <= 20'h398c6; 
			12'd136 : q <= 20'h98423; 
			12'd137 : q <= 20'h1b443; 
			12'd138 : q <= 20'h4110c; 
			12'd139 : q <= 20'h288c3; 
			12'd140 : q <= 20'h3052a; 
			12'd141 : q <= 20'h010cc; 
			12'd142 : q <= 20'h7b443; 
			12'd143 : q <= 20'h3b8a3; 
			12'd144 : q <= 20'h7b463; 
			12'd145 : q <= 20'h33903; 
			12'd146 : q <= 20'h7b463; 
			12'd147 : q <= 20'h13463; 
			12'd148 : q <= 20'h21d8c; 
			12'd149 : q <= 20'h49c46; 
			12'd150 : q <= 20'h424a2; 
			12'd151 : q <= 20'h41864; 
			12'd152 : q <= 20'h49848; 
			12'd153 : q <= 20'h39c66; 
			12'd154 : q <= 20'h58c63; 
			12'd155 : q <= 20'h290c1; 
			12'd156 : q <= 20'h29943; 
			12'd157 : q <= 20'h38cc9; 
			12'd158 : q <= 20'h31d21; 
			12'd159 : q <= 20'h12208; 
			12'd160 : q <= 20'h71846; 
			12'd161 : q <= 20'h094cf; 
			12'd162 : q <= 20'h500c9; 
			12'd163 : q <= 20'h318ee; 
			12'd164 : q <= 20'h69c66; 
			12'd165 : q <= 20'h0a1e4; 
			12'd166 : q <= 20'h5886a; 
			12'd167 : q <= 20'h19c86; 
			12'd168 : q <= 20'h68cca; 
			12'd169 : q <= 20'h29d0a; 
			12'd170 : q <= 20'h2118c; 
			12'd171 : q <= 20'h090c9; 
			12'd172 : q <= 20'h58c45; 
			12'd173 : q <= 20'h38c45; 
			12'd174 : q <= 20'h53843; 
			12'd175 : q <= 20'h2b0c2; 
			12'd176 : q <= 20'h4b843; 
			12'd177 : q <= 20'h22d86; 
			12'd178 : q <= 20'h5aca9; 
			12'd179 : q <= 20'h33c62; 
			12'd180 : q <= 20'h58065; 
			12'd181 : q <= 20'h294c7; 
			12'd182 : q <= 20'h68029; 
			12'd183 : q <= 20'h18888; 
			12'd184 : q <= 20'h6b086; 
			12'd185 : q <= 20'h1b086; 
			12'd186 : q <= 20'h6ac64; 
			12'd187 : q <= 20'h21083; 
			12'd188 : q <= 20'h39568; 
			12'd189 : q <= 20'h3a064; 
			12'd190 : q <= 20'h484c1; 
			12'd191 : q <= 20'h29463; 
			12'd192 : q <= 20'h02686; 
			12'd193 : q <= 20'h41865; 
			12'd194 : q <= 20'h58023; 
			12'd195 : q <= 20'h20882; 
			12'd196 : q <= 20'h61883; 
			12'd197 : q <= 20'h280c4; 
			12'd198 : q <= 20'h49c68; 
			12'd199 : q <= 20'h49c42; 
			12'd200 : q <= 20'h31dc4; 
			12'd201 : q <= 20'h01466; 
			12'd202 : q <= 20'h6ac64; 
			12'd203 : q <= 20'h22c64; 
			12'd204 : q <= 20'h2a588; 
			12'd205 : q <= 20'h4b023; 
			12'd206 : q <= 20'h53c44; 
			12'd207 : q <= 20'h39cc1; 
			12'd208 : q <= 20'h60cc6; 
			12'd209 : q <= 20'h01146; 
			12'd210 : q <= 20'h40d0e; 
			12'd211 : q <= 20'h210ef; 
			12'd212 : q <= 20'h608c8; 
			12'd213 : q <= 20'h108c8; 
			12'd214 : q <= 20'h13647; 
			12'd215 : q <= 20'h20d0e; 
			12'd216 : q <= 20'h90446; 
			12'd217 : q <= 20'h4ac43; 
			12'd218 : q <= 20'h90446; 
			12'd219 : q <= 20'h00446; 
			12'd220 : q <= 20'h09646; 
			12'd221 : q <= 20'h008c7; 
			12'd222 : q <= 20'h38cce; 
			12'd223 : q <= 20'h19daa; 
			12'd224 : q <= 20'h5bc42; 
			12'd225 : q <= 20'h12e04; 
			12'd226 : q <= 20'h69cc4; 
			12'd227 : q <= 20'h32869; 
			12'd228 : q <= 20'h71826; 
			12'd229 : q <= 20'h2a881; 
			12'd230 : q <= 20'h1a1e5; 
			12'd231 : q <= 20'h098a4; 
			12'd232 : q <= 20'h18626; 
			12'd233 : q <= 20'h31d02; 
			12'd234 : q <= 20'h49c62; 
			12'd235 : q <= 20'h41c62; 
			12'd236 : q <= 20'h42482; 
			12'd237 : q <= 20'h42083; 
			12'd238 : q <= 20'h494c4; 
			12'd239 : q <= 20'h43483; 
			12'd240 : q <= 20'h21d86; 
			12'd241 : q <= 20'h43883; 
			12'd242 : q <= 20'h49c63; 
			12'd243 : q <= 20'h39068; 
			12'd244 : q <= 20'h50066; 
			12'd245 : q <= 20'h30c88; 
			12'd246 : q <= 20'h70ccd; 
			12'd247 : q <= 20'h43466; 
			12'd248 : q <= 20'h70ccd; 
			12'd249 : q <= 20'h01d44; 
			12'd250 : q <= 20'h70ccd; 
			12'd251 : q <= 20'h00ccd; 
			12'd252 : q <= 20'h48481; 
			12'd253 : q <= 20'h40041; 
			12'd254 : q <= 20'h54084; 
			12'd255 : q <= 20'h49843; 
			12'd256 : q <= 20'h21582; 
			12'd257 : q <= 20'h41c65; 
			12'd258 : q <= 20'h31106; 
			12'd259 : q <= 20'h4944c; 
			12'd260 : q <= 20'h218c8; 
			12'd261 : q <= 20'h60905; 
			12'd262 : q <= 20'h02243; 
			12'd263 : q <= 20'h43088; 
			12'd264 : q <= 20'h00905; 
			12'd265 : q <= 20'h6ac64; 
			12'd266 : q <= 20'h2acc1; 
			12'd267 : q <= 20'h58c61; 
			12'd268 : q <= 20'h3b4a3; 
			12'd269 : q <= 20'h5ace6; 
			12'd270 : q <= 20'h12ce6; 
			12'd271 : q <= 20'h63846; 
			12'd272 : q <= 20'h43863; 
			12'd273 : q <= 20'h58065; 
			12'd274 : q <= 20'h30489; 
			12'd275 : q <= 20'h50cc1; 
			12'd276 : q <= 20'h42064; 
			12'd277 : q <= 20'h43082; 
			12'd278 : q <= 20'h2c882; 
			12'd279 : q <= 20'h10646; 
			12'd280 : q <= 20'h30062; 
			12'd281 : q <= 20'h6a0c2; 
			12'd282 : q <= 20'h32866; 
			12'd283 : q <= 20'h03684; 
			12'd284 : q <= 20'h39cc5; 
			12'd285 : q <= 20'h58042; 
			12'd286 : q <= 20'h0a0c2; 
			12'd287 : q <= 20'h00a82; 
			12'd288 : q <= 20'h3b8a3; 
			12'd289 : q <= 20'h3b4c6; 
			12'd290 : q <= 20'h4b043; 
			12'd291 : q <= 20'h82c26; 
			12'd292 : q <= 20'h1ac26; 
			12'd293 : q <= 20'h211cc; 
			12'd294 : q <= 20'h29063; 
			12'd295 : q <= 20'h60c63; 
			12'd296 : q <= 20'h31903; 
			12'd297 : q <= 20'h60c63; 
			12'd298 : q <= 20'h1848a; 
			12'd299 : q <= 20'h29d42; 
			12'd300 : q <= 20'h41c63; 
			12'd301 : q <= 20'h7b043; 
			12'd302 : q <= 20'h3a064; 
			12'd303 : q <= 20'h6902c; 
			12'd304 : q <= 20'h2158c; 
			12'd305 : q <= 20'h3b8e3; 
			12'd306 : q <= 20'h1b043; 
			12'd307 : q <= 20'h189c2; 
			12'd308 : q <= 20'h0046a; 
			12'd309 : q <= 20'h480c5; 
			12'd310 : q <= 20'h29cc2; 
			12'd311 : q <= 20'h384ca; 
			12'd312 : q <= 20'h08643; 
			12'd313 : q <= 20'h80c66; 
			12'd314 : q <= 20'h30ce6; 
			12'd315 : q <= 20'h21d82; 
			12'd316 : q <= 20'h0122a; 
			12'd317 : q <= 20'h191f0; 
			12'd318 : q <= 20'h3bcc4; 
			12'd319 : q <= 20'h78889; 
			12'd320 : q <= 20'h10c62; 
			12'd321 : q <= 20'h698e9; 
			12'd322 : q <= 20'h42c83; 
			12'd323 : q <= 20'h00a86; 
			12'd324 : q <= 20'h188ca; 
			12'd325 : q <= 20'h6a864; 
			12'd326 : q <= 20'h22864; 
			12'd327 : q <= 20'h394c3; 
			12'd328 : q <= 20'h398c8; 
			12'd329 : q <= 20'h02e86; 
			12'd330 : q <= 20'h23486; 
			12'd331 : q <= 20'h3010c; 
			12'd332 : q <= 20'h101e2; 
			12'd333 : q <= 20'h4b043; 
			12'd334 : q <= 20'h1b022; 
			12'd335 : q <= 20'h4ac43; 
			12'd336 : q <= 20'h38c61; 
			12'd337 : q <= 20'h89c66; 
			12'd338 : q <= 20'h38862; 
			12'd339 : q <= 20'h590a3; 
			12'd340 : q <= 20'h210a3; 
			12'd341 : q <= 20'h98c22; 
			12'd342 : q <= 20'h29483; 
			12'd343 : q <= 20'h89c66; 
			12'd344 : q <= 20'h01c66; 
			12'd345 : q <= 20'h708c9; 
			12'd346 : q <= 20'h010a6; 
			12'd347 : q <= 20'h514c2; 
			12'd348 : q <= 20'h214c2; 
			12'd349 : q <= 20'h40486; 
			12'd350 : q <= 20'h00866; 
			12'd351 : q <= 20'h31903; 
			12'd352 : q <= 20'h004a9; 
			12'd353 : q <= 20'h8008f; 
			12'd354 : q <= 20'h0a862; 
			12'd355 : q <= 20'h7102a; 
			12'd356 : q <= 20'h0048c; 
			12'd357 : q <= 20'h5ac82; 
			12'd358 : q <= 20'h2ac82; 
			12'd359 : q <= 20'h1a1e5; 
			12'd360 : q <= 20'h000ca; 
			12'd361 : q <= 20'h59062; 
			12'd362 : q <= 20'h43068; 
			12'd363 : q <= 20'h438a3; 
			12'd364 : q <= 20'h3b883; 
			12'd365 : q <= 20'h59062; 
			12'd366 : q <= 20'h1bdc4; 
			12'd367 : q <= 20'h10a04; 
			12'd368 : q <= 20'h020cc; 
			12'd369 : q <= 20'h29d42; 
			12'd370 : q <= 20'h49c45; 
			12'd371 : q <= 20'h69cc4; 
			12'd372 : q <= 20'h03502; 
			12'd373 : q <= 20'h69cc4; 
			12'd374 : q <= 20'h09cc4; 
			12'd375 : q <= 20'h6182c; 
			12'd376 : q <= 20'h49446; 
			12'd377 : q <= 20'h73043; 
			12'd378 : q <= 20'h23043; 
			12'd379 : q <= 20'h43083; 
			12'd380 : q <= 20'h28844; 
			12'd381 : q <= 20'h29563; 
			12'd382 : q <= 20'h3988c; 
			12'd383 : q <= 20'h63505; 
			12'd384 : q <= 20'h3982c; 
			12'd385 : q <= 20'h088c3; 
			12'd386 : q <= 20'h494ca; 
			12'd387 : q <= 20'h2950c; 
			12'd388 : q <= 20'h01e86; 
			12'd389 : q <= 20'h20842; 
			12'd390 : q <= 20'h24982; 
			12'd391 : q <= 20'h39090; 
			12'd392 : q <= 20'h398e8; 
			12'd393 : q <= 20'h30c61; 
			12'd394 : q <= 20'h5bc44; 
			12'd395 : q <= 20'h19488; 
			12'd396 : q <= 20'h384cc; 
			12'd397 : q <= 20'h218c2; 
			12'd398 : q <= 20'h81086; 
			12'd399 : q <= 20'h18ca2; 
			12'd400 : q <= 20'h4ac43; 
			12'd401 : q <= 20'h14082; 
			12'd402 : q <= 20'h3b4c6; 
			12'd403 : q <= 20'h38064; 
			12'd404 : q <= 20'h43c83; 
			12'd405 : q <= 20'h01086; 
			12'd406 : q <= 20'h29983; 
			12'd407 : q <= 20'h398ce; 
			12'd408 : q <= 20'h49c63; 
			12'd409 : q <= 20'h33044; 
			12'd410 : q <= 20'h530e6; 
			12'd411 : q <= 20'h081e2; 
			12'd412 : q <= 20'h700c6; 
			12'd413 : q <= 20'h28c61; 
			12'd414 : q <= 20'h700c6; 
			12'd415 : q <= 20'h00e8a; 
			12'd416 : q <= 20'h700c6; 
			12'd417 : q <= 20'h000c6; 
			12'd418 : q <= 20'h9bc22; 
			12'd419 : q <= 20'h00888; 
			12'd420 : q <= 20'h10644; 
			12'd421 : q <= 20'h43022; 
			12'd422 : q <= 20'h28946; 
			12'd423 : q <= 20'h49c44; 
			12'd424 : q <= 20'h49c63; 
			12'd425 : q <= 20'h21588; 
			12'd426 : q <= 20'h7bc83; 
			12'd427 : q <= 20'h44861; 
			12'd428 : q <= 20'h4b483; 
			12'd429 : q <= 20'h3b483; 
			12'd430 : q <= 20'h9bc22; 
			12'd431 : q <= 20'h03d04; 
			12'd432 : q <= 20'h48cc4; 
			12'd433 : q <= 20'h43883; 
			12'd434 : q <= 20'h1b9c6; 
			12'd435 : q <= 20'h30cc6; 
			12'd436 : q <= 20'h2ad46; 
			12'd437 : q <= 20'h1a864; 
			12'd438 : q <= 20'h6a442; 
			12'd439 : q <= 20'h28cc4; 
			12'd440 : q <= 20'h49c63; 
			12'd441 : q <= 20'h13043; 
			12'd442 : q <= 20'h4a06c; 
			12'd443 : q <= 20'h1b886; 
			12'd444 : q <= 20'h83c42; 
			12'd445 : q <= 20'h13c42; 
			12'd446 : q <= 20'h43083; 
			12'd447 : q <= 20'h01e81; 
			12'd448 : q <= 20'h39903; 
			12'd449 : q <= 20'h29d02; 
			12'd450 : q <= 20'h49c65; 
			12'd451 : q <= 20'h41c65; 
			12'd452 : q <= 20'h58465; 
			12'd453 : q <= 20'h30866; 
			12'd454 : q <= 20'h738c5; 
			12'd455 : q <= 20'h4a042; 
			12'd456 : q <= 20'h51c23; 
			12'd457 : q <= 20'h31842; 
			12'd458 : q <= 20'h12e44; 
			12'd459 : q <= 20'h31842; 
			12'd460 : q <= 20'h03e82; 
			12'd461 : q <= 20'h23843; 
			12'd462 : q <= 20'h43883; 
			12'd463 : q <= 20'h41c43; 
			12'd464 : q <= 20'h4a843; 
			12'd465 : q <= 20'h29144; 
			12'd466 : q <= 20'h49cc4; 
			12'd467 : q <= 20'h21c66; 
			12'd468 : q <= 20'h5bc84; 
			12'd469 : q <= 20'h3a082; 
			12'd470 : q <= 20'h68483; 
			12'd471 : q <= 20'h2bc84; 
			12'd472 : q <= 20'h49487; 
			12'd473 : q <= 20'h29903; 
			12'd474 : q <= 20'h4a442; 
			12'd475 : q <= 20'h3bca3; 
			12'd476 : q <= 20'h5a883; 
			12'd477 : q <= 20'h3250a; 
			12'd478 : q <= 20'h52cc2; 
			12'd479 : q <= 20'h22cc2; 
			12'd480 : q <= 20'h58d01; 
			12'd481 : q <= 20'h30c62; 
			12'd482 : q <= 20'h714c5; 
			12'd483 : q <= 20'h3944c; 
			12'd484 : q <= 20'h42c83; 
			12'd485 : q <= 20'h20443; 
			12'd486 : q <= 20'h90c46; 
			12'd487 : q <= 20'h00c46; 
			12'd488 : q <= 20'h4b043; 
			12'd489 : q <= 20'h3b483; 
			12'd490 : q <= 20'h90046; 
			12'd491 : q <= 20'h00046; 
			12'd492 : q <= 20'h438c3; 
			12'd493 : q <= 20'h39044; 
			12'd494 : q <= 20'h41486; 
			12'd495 : q <= 20'h31042; 
			12'd496 : q <= 20'h1b9c4; 
			12'd497 : q <= 20'h33cc2; 
			12'd498 : q <= 20'h73cc2; 
			12'd499 : q <= 20'h13188; 
			12'd500 : q <= 20'h39ce2; 
			12'd501 : q <= 20'h00a42; 
			12'd502 : q <= 20'h49845; 
			12'd503 : q <= 20'h39468; 
			12'd504 : q <= 20'h49864; 
			12'd505 : q <= 20'h23462; 
			12'd506 : q <= 20'h490c3; 
			12'd507 : q <= 20'h290c3; 
			12'd508 : q <= 20'h72ca2; 
			12'd509 : q <= 20'h088c9; 
			12'd510 : q <= 20'h718cd; 
			12'd511 : q <= 20'h199c8; 
			12'd512 : q <= 20'h8008b; 
			12'd513 : q <= 20'h1918c; 
			12'd514 : q <= 20'h590a3; 
			12'd515 : q <= 20'h22c82; 
			12'd516 : q <= 20'h51c42; 
			12'd517 : q <= 20'h41c42; 
			12'd518 : q <= 20'h4c462; 
			12'd519 : q <= 20'h29863; 
			12'd520 : q <= 20'h50063; 
			12'd521 : q <= 20'h298c2; 
			12'd522 : q <= 20'h64083; 
			12'd523 : q <= 20'h1b062; 
			12'd524 : q <= 20'h4b062; 
			12'd525 : q <= 20'h0ae04; 
			12'd526 : q <= 20'h61063; 
			12'd527 : q <= 20'h210a3; 
			12'd528 : q <= 20'h64083; 
			12'd529 : q <= 20'h29063; 
			12'd530 : q <= 20'h48042; 
			12'd531 : q <= 20'h42482; 
			12'd532 : q <= 20'h42083; 
			12'd533 : q <= 20'h034c3; 
			12'd534 : q <= 20'h83862; 
			12'd535 : q <= 20'h0ca42; 
			12'd536 : q <= 20'h83862; 
			12'd537 : q <= 20'h0b862; 
			12'd538 : q <= 20'h3b8c3; 
			12'd539 : q <= 20'h2b903; 
			12'd540 : q <= 20'h5188e; 
			12'd541 : q <= 20'h3188e; 
			12'd542 : q <= 20'h69443; 
			12'd543 : q <= 20'h3c0c1; 
			12'd544 : q <= 20'h4b063; 
			12'd545 : q <= 20'h38063; 
			12'd546 : q <= 20'h20212; 
			12'd547 : q <= 20'h0860e; 
			12'd548 : q <= 20'h1a5e4; 
			12'd549 : q <= 20'h330e3; 
			12'd550 : q <= 20'h73c43; 
			12'd551 : q <= 20'h10e0e; 
			12'd552 : q <= 20'h80892; 
			12'd553 : q <= 20'h23c43; 
			12'd554 : q <= 20'h80892; 
			12'd555 : q <= 20'h08503; 
			12'd556 : q <= 20'h42c83; 
			12'd557 : q <= 20'h2aca9; 
			12'd558 : q <= 20'h8008b; 
			12'd559 : q <= 20'h380c1; 
			12'd560 : q <= 20'h80c67; 
			12'd561 : q <= 20'h08c67; 
			12'd562 : q <= 20'h3a0cc; 
			12'd563 : q <= 20'h0008b; 
			12'd564 : q <= 20'h700d4; 
			12'd565 : q <= 20'h00c22; 
			12'd566 : q <= 20'h29548; 
			12'd567 : q <= 20'h21d84; 
			12'd568 : q <= 20'h104c4; 
			12'd569 : q <= 20'h49cc4; 
			12'd570 : q <= 20'h29846; 
			12'd571 : q <= 20'h4c0c4; 
			12'd572 : q <= 20'h4904c; 
			12'd573 : q <= 20'h384d2; 
			12'd574 : q <= 20'h23182; 
			12'd575 : q <= 20'h420c2; 
			12'd576 : q <= 20'h40066; 
			12'd577 : q <= 20'h5c862; 
			12'd578 : q <= 20'h08624; 
			12'd579 : q <= 20'h5a08c; 
			12'd580 : q <= 20'h43883; 
			12'd581 : q <= 20'h60c51; 
			12'd582 : q <= 20'h21cc1; 
			12'd583 : q <= 20'h90c43; 
			12'd584 : q <= 20'h41064; 
			12'd585 : q <= 20'h2158a; 
			12'd586 : q <= 20'h2c882; 
			12'd587 : q <= 20'h88866; 
			12'd588 : q <= 20'h39cc6; 
			12'd589 : q <= 20'h88866; 
			12'd590 : q <= 20'h40064; 
			12'd591 : q <= 20'h4b843; 
			12'd592 : q <= 20'h030c3; 
			12'd593 : q <= 20'h43883; 
			12'd594 : q <= 20'h1b043; 
			12'd595 : q <= 20'h29987; 
			12'd596 : q <= 20'h00866; 
			12'd597 : q <= 20'h71823; 
			12'd598 : q <= 20'h1006e; 
			12'd599 : q <= 20'h638a6; 
			12'd600 : q <= 20'h238a6; 
			12'd601 : q <= 20'h5a842; 
			12'd602 : q <= 20'h2806e; 
			12'd603 : q <= 20'h53c43; 
			12'd604 : q <= 20'h00843; 
			12'd605 : q <= 20'h2ad86; 
			12'd606 : q <= 20'h32c69; 
			12'd607 : q <= 20'h5a842; 
			12'd608 : q <= 20'h29823; 
			12'd609 : q <= 20'h225a3; 
			12'd610 : q <= 20'h09de6; 
			12'd611 : q <= 20'h21586; 
			12'd612 : q <= 20'h42883; 
			12'd613 : q <= 20'h7b823; 
			12'd614 : q <= 20'h0aca3; 
			12'd615 : q <= 20'h384ec; 
			12'd616 : q <= 20'h004ca; 
			12'd617 : q <= 20'h80483; 
			12'd618 : q <= 20'h29443; 
			12'd619 : q <= 20'h60865; 
			12'd620 : q <= 20'h00c86; 
			12'd621 : q <= 20'h43082; 
			12'd622 : q <= 20'h44861; 
			12'd623 : q <= 20'h5a842; 
			12'd624 : q <= 20'h3a842; 
			12'd625 : q <= 20'h5ac84; 
			12'd626 : q <= 20'h43068; 
			12'd627 : q <= 20'h680c3; 
			12'd628 : q <= 20'h42064; 
			12'd629 : q <= 20'h29d4a; 
			12'd630 : q <= 20'h1c902; 
			12'd631 : q <= 20'h508c8; 
			12'd632 : q <= 20'h208c8; 
			12'd633 : q <= 20'h58067; 
			12'd634 : q <= 20'h3ac41; 
			12'd635 : q <= 20'h7b823; 
			12'd636 : q <= 20'h3bc42; 
			12'd637 : q <= 20'h7b823; 
			12'd638 : q <= 20'h30067; 
			12'd639 : q <= 20'h90447; 
			12'd640 : q <= 20'h10114; 
			12'd641 : q <= 20'h181e6; 
			12'd642 : q <= 20'h20d82; 
			12'd643 : q <= 20'h80085; 
			12'd644 : q <= 20'h38064; 
			12'd645 : q <= 20'h80085; 
			12'd646 : q <= 20'h09ccd; 
			12'd647 : q <= 20'h80085; 
			12'd648 : q <= 20'h00085; 
			12'd649 : q <= 20'h73066; 
			12'd650 : q <= 20'h1b066; 
			12'd651 : q <= 20'h80483; 
			12'd652 : q <= 20'h41c4a; 
			12'd653 : q <= 20'h5ac84; 
			12'd654 : q <= 20'h00483; 
			12'd655 : q <= 20'h69023; 
			12'd656 : q <= 20'h3bc65; 
			12'd657 : q <= 20'h49c65; 
			12'd658 : q <= 20'h41c65; 
			12'd659 : q <= 20'h5188e; 
			12'd660 : q <= 20'h014a6; 
			12'd661 : q <= 20'h494c4; 
			12'd662 : q <= 20'h0024a; 
			12'd663 : q <= 20'h5188e; 
			12'd664 : q <= 20'h3188e; 
			12'd665 : q <= 20'h69023; 
			12'd666 : q <= 20'h28443; 
			12'd667 : q <= 20'h90452; 
			12'd668 : q <= 20'h10483; 
			12'd669 : q <= 20'h90452; 
			12'd670 : q <= 20'h0b886; 
			12'd671 : q <= 20'h52ce6; 
			12'd672 : q <= 20'h028ca; 
			12'd673 : q <= 20'h58064; 
			12'd674 : q <= 20'h2a8a6; 
			12'd675 : q <= 20'h71828; 
			12'd676 : q <= 20'h09e46; 
			12'd677 : q <= 20'h49c42; 
			12'd678 : q <= 20'h2a485; 
			12'd679 : q <= 20'h398c3; 
			12'd680 : q <= 20'h08244; 
			12'd681 : q <= 20'h3bc44; 
			12'd682 : q <= 20'h08269; 
			12'd683 : q <= 20'h19c66; 
			12'd684 : q <= 20'h69c84; 
			12'd685 : q <= 20'h19c84; 
			12'd686 : q <= 20'h49948; 
			12'd687 : q <= 20'h1a1cc; 
			12'd688 : q <= 20'h3154c; 
			12'd689 : q <= 20'h4ac43; 
			12'd690 : q <= 20'h494c5; 
			12'd691 : q <= 20'h49044; 
			12'd692 : q <= 20'h494c5; 
			12'd693 : q <= 20'h294c5; 
			12'd694 : q <= 20'h588c1; 
			12'd695 : q <= 20'h188c1; 
			12'd696 : q <= 20'h69443; 
			12'd697 : q <= 20'h02824; 
			12'd698 : q <= 20'h69443; 
			12'd699 : q <= 20'h44862; 
			12'd700 : q <= 20'h33d22; 
			12'd701 : q <= 20'h43883; 
			12'd702 : q <= 20'h91044; 
			12'd703 : q <= 20'h29443; 
			12'd704 : q <= 20'h7c062; 
			12'd705 : q <= 20'h00069; 
			12'd706 : q <= 20'h49c63; 
			12'd707 : q <= 20'h41c63; 
			12'd708 : q <= 20'h49446; 
			12'd709 : q <= 20'h41864; 
			12'd710 : q <= 20'h3990c; 
			12'd711 : q <= 20'h2990c; 
			12'd712 : q <= 20'h61063; 
			12'd713 : q <= 20'h14062; 
			12'd714 : q <= 20'h61063; 
			12'd715 : q <= 20'h130c6; 
			12'd716 : q <= 20'h3b4c3; 
			12'd717 : q <= 20'h338c3; 
			12'd718 : q <= 20'h73ca3; 
			12'd719 : q <= 20'h29063; 
			12'd720 : q <= 20'h73ca3; 
			12'd721 : q <= 20'h28cc2; 
			12'd722 : q <= 20'h43c83; 
			12'd723 : q <= 20'h0bca3; 
			12'd724 : q <= 20'h43486; 
			12'd725 : q <= 20'h3a063; 
			12'd726 : q <= 20'h600a4; 
			12'd727 : q <= 20'h00a82; 
			12'd728 : q <= 20'h08244; 
			12'd729 : q <= 20'h20cc1; 
			12'd730 : q <= 20'h249a2; 
			12'd731 : q <= 20'h12866; 
			12'd732 : q <= 20'h730c8; 
			12'd733 : q <= 20'h23546; 
			12'd734 : q <= 20'h73022; 
			12'd735 : q <= 20'h43483; 
			12'd736 : q <= 20'h73042; 
			12'd737 : q <= 20'h23042; 
			12'd738 : q <= 20'h43122; 
			12'd739 : q <= 20'h4b843; 
			12'd740 : q <= 20'h5a866; 
			12'd741 : q <= 20'h2992c; 
			12'd742 : q <= 20'h5a866; 
			12'd743 : q <= 20'h32866; 
			12'd744 : q <= 20'h29163; 
			12'd745 : q <= 20'h384aa; 
			12'd746 : q <= 20'h12242; 
			12'd747 : q <= 20'h3c4a3; 
			12'd748 : q <= 20'h2a581; 
			12'd749 : q <= 20'h038c6; 
			12'd750 : q <= 20'h2a581; 
			12'd751 : q <= 20'h1a581; 
			12'd752 : q <= 20'h728c7; 
			12'd753 : q <= 20'h08202; 
			12'd754 : q <= 20'h52549; 
			12'd755 : q <= 20'h00542; 
			12'd756 : q <= 20'h88c43; 
			12'd757 : q <= 20'h08c43; 
			12'd758 : q <= 20'h49c66; 
			12'd759 : q <= 20'h31483; 
			12'd760 : q <= 20'h394c6; 
			12'd761 : q <= 20'h1918c; 
			12'd762 : q <= 20'h488cf; 
			12'd763 : q <= 20'h108d1; 
			12'd764 : q <= 20'h728c7; 
			12'd765 : q <= 20'h028c7; 
			12'd766 : q <= 20'h488cf; 
			12'd767 : q <= 20'h288cf; 
			12'd768 : q <= 20'h8a466; 
			12'd769 : q <= 20'h31cc6; 
			12'd770 : q <= 20'h0aa46; 
			12'd771 : q <= 20'h02549; 
			12'd772 : q <= 20'h43c83; 
			12'd773 : q <= 20'h2b064; 
			12'd774 : q <= 20'h18e0c; 
			12'd775 : q <= 20'h0858c; 
			12'd776 : q <= 20'h51044; 
			12'd777 : q <= 20'h02542; 
			12'd778 : q <= 20'h4ac63; 
			12'd779 : q <= 20'h1b122; 
			12'd780 : q <= 20'h4a442; 
			12'd781 : q <= 20'h191a6; 
			12'd782 : q <= 20'h49cc4; 
			12'd783 : q <= 20'h080c8; 
			12'd784 : q <= 20'h4944c; 
			12'd785 : q <= 20'h2106a; 
			12'd786 : q <= 20'h34503; 
			12'd787 : q <= 20'h01546; 
			12'd788 : q <= 20'h68862; 
			12'd789 : q <= 20'h39485; 
			12'd790 : q <= 20'h63866; 
			12'd791 : q <= 20'h0ad02; 
			12'd792 : q <= 20'h3b4c3; 
			12'd793 : q <= 20'h01466; 
			12'd794 : q <= 20'h68862; 
			12'd795 : q <= 20'h23886; 
			12'd796 : q <= 20'h68862; 
			12'd797 : q <= 20'h4088c; 
			12'd798 : q <= 20'h700c8; 
			12'd799 : q <= 20'h3c462; 
			12'd800 : q <= 20'h43082; 
			12'd801 : q <= 20'h3010c; 
			12'd802 : q <= 20'h7004a; 
			12'd803 : q <= 20'h28d06; 
			12'd804 : q <= 20'h700ca; 
			12'd805 : q <= 20'h4b822; 
			12'd806 : q <= 20'h7a883; 
			12'd807 : q <= 20'h43843; 
			12'd808 : q <= 20'h1b5c4; 
			12'd809 : q <= 20'h0a883; 
			12'd810 : q <= 20'h4acc1; 
			12'd811 : q <= 20'h2acc1; 
			12'd812 : q <= 20'h1960f; 
			12'd813 : q <= 20'h33082; 
			12'd814 : q <= 20'h2118a; 
			12'd815 : q <= 20'h41864; 
			12'd816 : q <= 20'h43088; 
			12'd817 : q <= 20'h43883; 
			12'd818 : q <= 20'h60862; 
			12'd819 : q <= 20'h43c62; 
			12'd820 : q <= 20'h3012e; 
			12'd821 : q <= 20'h49843; 
			12'd822 : q <= 20'h52043; 
			12'd823 : q <= 20'h02486; 
			12'd824 : q <= 20'h30102; 
			12'd825 : q <= 20'h338e3; 
			12'd826 : q <= 20'h42909; 
			12'd827 : q <= 20'h28862; 
			12'd828 : q <= 20'h704c8; 
			12'd829 : q <= 20'h004c8; 
			12'd830 : q <= 20'h08a46; 
			12'd831 : q <= 20'h48c41; 
			12'd832 : q <= 20'h68886; 
			12'd833 : q <= 20'h29063; 
			12'd834 : q <= 20'h69423; 
			12'd835 : q <= 20'h140a3; 
			12'd836 : q <= 20'h68886; 
			12'd837 : q <= 20'h18886; 
			12'd838 : q <= 20'h69422; 
			12'd839 : q <= 20'h29442; 
			12'd840 : q <= 20'h6a442; 
			12'd841 : q <= 20'h2a442; 
			12'd842 : q <= 20'h6c462; 
			12'd843 : q <= 20'h34084; 
			12'd844 : q <= 20'h4c043; 
			12'd845 : q <= 20'h03526; 
			12'd846 : q <= 20'h4b846; 
			12'd847 : q <= 20'h4bc43; 
			12'd848 : q <= 20'h0aa46; 
			12'd849 : q <= 20'h42c82; 
			12'd850 : q <= 20'h3a4c2; 
			12'd851 : q <= 20'h42043; 
			12'd852 : q <= 20'h89464; 
			12'd853 : q <= 20'h0ce41; 
			12'd854 : q <= 20'h48062; 
			12'd855 : q <= 20'h0a026; 
			12'd856 : q <= 20'h64503; 
			12'd857 : q <= 20'h01464; 
			12'd858 : q <= 20'h49c43; 
			12'd859 : q <= 20'h3ac42; 
			12'd860 : q <= 20'h58c45; 
			12'd861 : q <= 20'h38c45; 
			12'd862 : q <= 20'h7b443; 
			12'd863 : q <= 20'h29843; 
			12'd864 : q <= 20'h24de1; 
			12'd865 : q <= 20'h0cde1; 
			12'd866 : q <= 20'h7b443; 
			12'd867 : q <= 20'h2808f; 
			12'd868 : q <= 20'h49845; 
			12'd869 : q <= 20'h49447; 
			12'd870 : q <= 20'h82c63; 
			12'd871 : q <= 20'h0ac63; 
			12'd872 : q <= 20'h31903; 
			12'd873 : q <= 20'h03cc2; 
			12'd874 : q <= 20'h08246; 
			12'd875 : q <= 20'h30064; 
			12'd876 : q <= 20'h7288a; 
			12'd877 : q <= 20'h18862; 
			12'd878 : q <= 20'h58842; 
			12'd879 : q <= 20'h1288a; 
			12'd880 : q <= 20'h03686; 
			12'd881 : q <= 20'h0144f; 
			12'd882 : q <= 20'h09e44; 
			12'd883 : q <= 20'h00051; 
			12'd884 : q <= 20'h11a06; 
			12'd885 : q <= 20'h43823; 
			12'd886 : q <= 20'h43c82; 
			12'd887 : q <= 20'h28902; 
			12'd888 : q <= 20'h32d06; 
			12'd889 : q <= 20'h4b442; 
			12'd890 : q <= 20'h91046; 
			12'd891 : q <= 20'h4b042; 
			12'd892 : q <= 20'h91046; 
			12'd893 : q <= 20'h4b423; 
			12'd894 : q <= 20'h91046; 
			12'd895 : q <= 20'h01046; 
			12'd896 : q <= 20'h4b063; 
			12'd897 : q <= 20'h1b443; 
			12'd898 : q <= 20'h6b483; 
			12'd899 : q <= 20'h29063; 
			12'd900 : q <= 20'h28946; 
			12'd901 : q <= 20'h1b483; 
			12'd902 : q <= 20'h19de5; 
			12'd903 : q <= 20'h19d82; 
			12'd904 : q <= 20'h50c69; 
			12'd905 : q <= 20'h41886; 
			12'd906 : q <= 20'h49c83; 
			12'd907 : q <= 20'h02489; 
			12'd908 : q <= 20'h4b465; 
			12'd909 : q <= 20'h39cc3; 
			12'd910 : q <= 20'h49c65; 
			12'd911 : q <= 20'h29d02; 
			12'd912 : q <= 20'h2a582; 
			12'd913 : q <= 20'h29943; 
			12'd914 : q <= 20'h53061; 
			12'd915 : q <= 20'h0056f; 
			12'd916 : q <= 20'h08246; 
			12'd917 : q <= 20'h39cc1; 
			12'd918 : q <= 20'h2c0c4; 
			12'd919 : q <= 20'h31528; 
			12'd920 : q <= 20'h2a846; 
			12'd921 : q <= 20'h3990a; 
			12'd922 : q <= 20'h2990a; 
			12'd923 : q <= 20'h49442; 
			12'd924 : q <= 20'h2b102; 
			12'd925 : q <= 20'h50902; 
			12'd926 : q <= 20'h2004a; 
			12'd927 : q <= 20'h4a842; 
			12'd928 : q <= 20'h121e3; 
			12'd929 : q <= 20'h43483; 
			12'd930 : q <= 20'h38862; 
			12'd931 : q <= 20'h3b4c3; 
			12'd932 : q <= 20'h4a442; 
			12'd933 : q <= 20'h88866; 
			12'd934 : q <= 20'h09464; 
			12'd935 : q <= 20'h72086; 
			12'd936 : q <= 20'h09068; 
			12'd937 : q <= 20'h43486; 
			12'd938 : q <= 20'h1b842; 
			12'd939 : q <= 20'h72086; 
			12'd940 : q <= 20'h12086; 
			12'd941 : q <= 20'h53826; 
			12'd942 : q <= 20'h39466; 
			12'd943 : q <= 20'h58846; 
			12'd944 : q <= 20'h318c5; 
			12'd945 : q <= 20'h88466; 
			12'd946 : q <= 20'h41c65; 
			12'd947 : q <= 20'h4c862; 
			12'd948 : q <= 20'h44862; 
			12'd949 : q <= 20'h60ca2; 
			12'd950 : q <= 20'h384ac; 
			12'd951 : q <= 20'h08244; 
			12'd952 : q <= 20'h20842; 
			12'd953 : q <= 20'h5b882; 
			12'd954 : q <= 20'h00866; 
			12'd955 : q <= 20'h49c43; 
			12'd956 : q <= 20'h29423; 
			12'd957 : q <= 20'h528c1; 
			12'd958 : q <= 20'h228c1; 
			12'd959 : q <= 20'h4c463; 
			12'd960 : q <= 20'h23823; 
			12'd961 : q <= 20'h61463; 
			12'd962 : q <= 20'h21583; 
			12'd963 : q <= 20'h4a043; 
			12'd964 : q <= 20'h22463; 
			12'd965 : q <= 20'h30131; 
			12'd966 : q <= 20'h4b023; 
			12'd967 : q <= 20'h4944f; 
			12'd968 : q <= 20'h43843; 
			12'd969 : q <= 20'h53823; 
			12'd970 : q <= 20'h384c5; 
			12'd971 : q <= 20'h00282; 
			12'd972 : q <= 20'h134a3; 
			12'd973 : q <= 20'h4ac43; 
			12'd974 : q <= 20'h1152f; 
			12'd975 : q <= 20'h2818a; 
			12'd976 : q <= 20'h28443; 
			12'd977 : q <= 20'h51cc1; 
			12'd978 : q <= 20'h1844a; 
			12'd979 : q <= 20'h69c41; 
			12'd980 : q <= 20'h23486; 
			12'd981 : q <= 20'h69c41; 
			12'd982 : q <= 20'h29c41; 
			12'd983 : q <= 20'h13244; 
			12'd984 : q <= 20'h29c42; 
			12'd985 : q <= 20'h80c82; 
			12'd986 : q <= 20'h00852; 
			12'd987 : q <= 20'h08a44; 
			12'd988 : q <= 20'h4b823; 
			12'd989 : q <= 20'h13244; 
			12'd990 : q <= 20'h03244; 
			12'd991 : q <= 20'h590a3; 
			12'd992 : q <= 20'h310e3; 
			12'd993 : q <= 20'h6c463; 
			12'd994 : q <= 20'h40464; 
			12'd995 : q <= 20'h59044; 
			12'd996 : q <= 20'h04523; 
			12'd997 : q <= 20'h58048; 
			12'd998 : q <= 20'h020cc; 
			12'd999 : q <= 20'h51c8c; 
			12'd1000 :q  <= 20'h28d0e; 
			12'd1001 :q  <= 20'h728c1; 
			12'd1002 :q  <= 20'h01144; 
			12'd1003 :q  <= 20'h500a8; 
			12'd1004 :q  <= 20'h40488; 
			12'd1005 :q  <= 20'h4acc1; 
			12'd1006 :q  <= 20'h42464; 
			12'd1007 :q  <= 20'h91046; 
			12'd1008 :q  <= 20'h42064; 
			12'd1009 :q  <= 20'h385a3; 
			12'd1010 :q  <= 20'h3b4c1; 
			12'd1011 :q  <= 20'h62c66; 
			12'd1012 :q  <= 20'h2acc1; 
			12'd1013 :q  <= 20'h0924a; 
			12'd1014 :q  <= 20'h41889; 
			12'd1015 :q  <= 20'h41883; 
			12'd1016 :q  <= 20'h41c63; 
			12'd1017 :q  <= 20'h73c83; 
			12'd1018 :q  <= 20'h2a86a; 
			12'd1019 :q  <= 20'h43c83; 
			12'd1020 :q  <= 20'h02026; 
			12'd1021 :q  <= 20'h53c23; 
			12'd1022 :q  <= 20'h13c83; 
			12'd1023 :q  <= 20'h90c48; 
			12'd1024 :q  <= 20'h00c48; 
			12'd1025 :q  <= 20'h19dca; 
			12'd1026 :q  <= 20'h01e63; 
			12'd1027 :q  <= 20'h61863; 
			12'd1028 :q  <= 20'h01823; 
			12'd1029 :q  <= 20'h61863; 
			12'd1030 :q  <= 20'h29863; 
			12'd1031 :q  <= 20'h40882; 
			12'd1032 :q  <= 20'h30c8c; 
			12'd1033 :q  <= 20'h69843; 
			12'd1034 :q  <= 20'h02a84; 
			12'd1035 :q  <= 20'h1022e; 
			12'd1036 :q  <= 20'h000ca; 
			12'd1037 :q  <= 20'h718c4; 
			12'd1038 :q  <= 20'h018c4; 
			12'd1039 :q  <= 20'h688e2; 
			12'd1040 :q  <= 20'h008e2; 
			12'd1041 :q  <= 20'h32dc2; 
			12'd1042 :q  <= 20'h41442; 
			12'd1043 :q  <= 20'h6a443; 
			12'd1044 :q  <= 20'h0846c; 
			12'd1045 :q  <= 20'h89023; 
			12'd1046 :q  <= 20'h11023; 
			12'd1047 :q  <= 20'h71423; 
			12'd1048 :q  <= 20'h3c043; 
			12'd1049 :q  <= 20'h43486; 
			12'd1050 :q  <= 20'h29423; 
			12'd1051 :q  <= 20'h80094; 
			12'd1052 :q  <= 20'h28446; 
			12'd1053 :q  <= 20'h29144; 
			12'd1054 :q  <= 20'h7888c; 
			12'd1055 :q  <= 20'h3988c; 
			12'd1056 :q  <= 20'h71428; 
			12'd1057 :q  <= 20'h091ca; 
			12'd1058 :q  <= 20'h598ce; 
			12'd1059 :q  <= 20'h198ce; 
			12'd1060 :q  <= 20'h225e2; 
			12'd1061 :q  <= 20'h3b8c3; 
			12'd1062 :q  <= 20'h30dc4; 
			12'd1063 :q  <= 20'h0a5e2; 
			12'd1064 :q  <= 20'h32d09; 
			12'd1065 :q  <= 20'h39068; 
			12'd1066 :q  <= 20'h71846; 
			12'd1067 :q  <= 20'h29cc4; 
			12'd1068 :q  <= 20'h08653; 
			12'd1069 :q  <= 20'h088c5; 
			12'd1070 :q  <= 20'h644c2; 
			12'd1071 :q  <= 20'h144c2; 
			12'd1072 :q  <= 20'h88c66; 
			12'd1073 :q  <= 20'h44463; 
			12'd1074 :q  <= 20'h53446; 
			12'd1075 :q  <= 20'h3b4c3; 
			12'd1076 :q  <= 20'h88c66; 
			12'd1077 :q  <= 20'h43443; 
			12'd1078 :q  <= 20'h48cc2; 
			12'd1079 :q  <= 20'h00c66; 
			12'd1080 :q  <= 20'h41486; 
			12'd1081 :q  <= 20'h29462; 
			12'd1082 :q  <= 20'h50464; 
			12'd1083 :q  <= 20'h088a9; 
			12'd1084 :q  <= 20'h69843; 
			12'd1085 :q  <= 20'h019c3; 
			12'd1086 :q  <= 20'h12e48; 
			12'd1087 :q  <= 20'h29843; 
			12'd1088 :q  <= 20'h51882; 
			12'd1089 :q  <= 20'h31882; 
			12'd1090 :q  <= 20'h50464; 
			12'd1091 :q  <= 20'h38447; 
			12'd1092 :q  <= 20'h209ee; 
			12'd1093 :q  <= 20'h41c62; 
			12'd1094 :q  <= 20'h10e44; 
			12'd1095 :q  <= 20'h49c42; 
			12'd1096 :q  <= 20'h6a443; 
			12'd1097 :q  <= 20'h288c2; 
			12'd1098 :q  <= 20'h49447; 
			12'd1099 :q  <= 20'h2a443; 
			12'd1100 :q  <= 20'h301d2; 
			12'd1101 :q  <= 20'h140c3; 
			12'd1102 :q  <= 20'h49c66; 
			12'd1103 :q  <= 20'h3a083; 
			12'd1104 :q  <= 20'h3b0c3; 
			12'd1105 :q  <= 20'h4b043; 
			12'd1106 :q  <= 20'h3b0c2; 
			12'd1107 :q  <= 20'h2ac86; 
			12'd1108 :q  <= 20'h5b0e2; 
			12'd1109 :q  <= 20'h32906; 
			12'd1110 :q  <= 20'h5a864; 
			12'd1111 :q  <= 20'h4c043; 
			12'd1112 :q  <= 20'h68c29; 
			12'd1113 :q  <= 20'h0b5c6; 
			12'd1114 :q  <= 20'h69826; 
			12'd1115 :q  <= 20'h01068; 
			12'd1116 :q  <= 20'h90052; 
			12'd1117 :q  <= 20'h10cc2; 
			12'd1118 :q  <= 20'h48106; 
			12'd1119 :q  <= 20'h31826; 
			12'd1120 :q  <= 20'h720c3; 
			12'd1121 :q  <= 20'h00052; 
			12'd1122 :q  <= 20'h0ca42; 
			12'd1123 :q  <= 20'h1bc42; 
			12'd1124 :q  <= 20'h438a3; 
			12'd1125 :q  <= 20'h43843; 
			12'd1126 :q  <= 20'h60c63; 
			12'd1127 :q  <= 20'h394c2; 
			12'd1128 :q  <= 20'h794a2; 
			12'd1129 :q  <= 20'h014a2; 
			12'd1130 :q  <= 20'h8b826; 
			12'd1131 :q  <= 20'h12523; 
			12'd1132 :q  <= 20'h60c63; 
			12'd1133 :q  <= 20'h00092; 
			12'd1134 :q  <= 20'h89823; 
			12'd1135 :q  <= 20'h13826; 
			12'd1136 :q  <= 20'h9a022; 
			12'd1137 :q  <= 20'h28c63; 
			12'd1138 :q  <= 20'h4c043; 
			12'd1139 :q  <= 20'h11823; 
			12'd1140 :q  <= 20'h61102; 
			12'd1141 :q  <= 20'h01102; 
			12'd1142 :q  <= 20'h14244; 
			12'd1143 :q  <= 20'h3bc44; 
			12'd1144 :q  <= 20'h201c3; 
			12'd1145 :q  <= 20'h00094; 
			12'd1146 :q  <= 20'h61088; 
			12'd1147 :q  <= 20'h31c42; 
			12'd1148 :q  <= 20'h51843; 
			12'd1149 :q  <= 20'h41c62; 
			12'd1150 :q  <= 20'h408cc; 
			12'd1151 :q  <= 20'h2016c; 
			12'd1152 :q  <= 20'h724cb; 
			12'd1153 :q  <= 20'h03883; 
			12'd1154 :q  <= 20'h4a843; 
			12'd1155 :q  <= 20'h2ac62; 
			12'd1156 :q  <= 20'h4bc63; 
			12'd1157 :q  <= 20'h42064; 
			12'd1158 :q  <= 20'h4bc63; 
			12'd1159 :q  <= 20'h39c62; 
			12'd1160 :q  <= 20'h12a04; 
			12'd1161 :q  <= 20'h10c91; 
			12'd1162 :q  <= 20'h7b447; 
			12'd1163 :q  <= 20'h108c1; 
			12'd1164 :q  <= 20'h28984; 
			12'd1165 :q  <= 20'h3010c; 
			12'd1166 :q  <= 20'h69c42; 
			12'd1167 :q  <= 20'h03286; 
			12'd1168 :q  <= 20'h71c43; 
			12'd1169 :q  <= 20'h0212c; 
			12'd1170 :q  <= 20'h18202; 
			12'd1171 :q  <= 20'h33c63; 
			12'd1172 :q  <= 20'h43cc3; 
			12'd1173 :q  <= 20'h02826; 
			12'd1174 :q  <= 20'h52483; 
			12'd1175 :q  <= 20'h4bc43; 
			12'd1176 :q  <= 20'h29d41; 
			12'd1177 :q  <= 20'h20193; 
			12'd1178 :q  <= 20'h01a86; 
			12'd1179 :q  <= 20'h19842; 
			12'd1180 :q  <= 20'h79842; 
			12'd1181 :q  <= 20'h19842; 
			12'd1182 :q  <= 20'h7102c; 
			12'd1183 :q  <= 20'h1160a; 
			12'd1184 :q  <= 20'h4c462; 
			12'd1185 :q  <= 20'h09042; 
			12'd1186 :q  <= 20'h281e5; 
			12'd1187 :q  <= 20'h001e5; 
			12'd1188 :q  <= 20'h58851; 
			12'd1189 :q  <= 20'h38851; 
			12'd1190 :q  <= 20'h7ac49; 
			12'd1191 :q  <= 20'h1ac49; 
			12'd1192 :q  <= 20'h2c1c4; 
			12'd1193 :q  <= 20'h09241; 
			12'd1194 :q  <= 20'h69cc4; 
			12'd1195 :q  <= 20'h4a04c; 
			12'd1196 :q  <= 20'h604c6; 
			12'd1197 :q  <= 20'h288c6; 
			12'd1198 :q  <= 20'h4c0c4; 
			12'd1199 :q  <= 20'h08a43; 
			12'd1200 :q  <= 20'h3912a; 
			12'd1201 :q  <= 20'h2a484; 
			12'd1202 :q  <= 20'h5a866; 
			12'd1203 :q  <= 20'h3aca3; 
			12'd1204 :q  <= 20'h3acc6; 
			12'd1205 :q  <= 20'h00149; 
			12'd1206 :q  <= 20'h6b826; 
			12'd1207 :q  <= 20'h00866; 
			12'd1208 :q  <= 20'h43883; 
			12'd1209 :q  <= 20'h33826; 
			12'd1210 :q  <= 20'h4bc43; 
			12'd1211 :q  <= 20'h31063; 
			12'd1212 :q  <= 20'h48163; 
			12'd1213 :q  <= 20'h01a83; 
			12'd1214 :q  <= 20'h50422; 
			12'd1215 :q  <= 20'h49846; 
			12'd1216 :q  <= 20'h2a181; 
			12'd1217 :q  <= 20'h1a181; 
			12'd1218 :q  <= 20'h49c65; 
			12'd1219 :q  <= 20'h1a4c2; 
			12'd1220 :q  <= 20'h62463; 
			12'd1221 :q  <= 20'h380c1; 
			12'd1222 :q  <= 20'h62463; 
			12'd1223 :q  <= 20'h3a841; 
			12'd1224 :q  <= 20'h3112d; 
			12'd1225 :q  <= 20'h32082; 
			12'd1226 :q  <= 20'h80886; 
			12'd1227 :q  <= 20'h044c3; 
			12'd1228 :q  <= 20'h5286a; 
			12'd1229 :q  <= 20'h41c65; 
			12'd1230 :q  <= 20'h51083; 
			12'd1231 :q  <= 20'h41068; 
			12'd1232 :q  <= 20'h3192d; 
			12'd1233 :q  <= 20'h3010c; 
			12'd1234 :q  <= 20'h708c8; 
			12'd1235 :q  <= 20'h30066; 
			12'd1236 :q  <= 20'h708c8; 
			12'd1237 :q  <= 20'h014c6; 
			12'd1238 :q  <= 20'h4b0c2; 
			12'd1239 :q  <= 20'h44462; 
			12'd1240 :q  <= 20'h59842; 
			12'd1241 :q  <= 20'h0a642; 
			12'd1242 :q  <= 20'h59842; 
			12'd1243 :q  <= 20'h19188; 
			12'd1244 :q  <= 20'h6aca3; 
			12'd1245 :q  <= 20'h4a843; 
			12'd1246 :q  <= 20'h71c43; 
			12'd1247 :q  <= 20'h29023; 
			12'd1248 :q  <= 20'h69043; 
			12'd1249 :q  <= 20'h29043; 
			12'd1250 :q  <= 20'h4a043; 
			12'd1251 :q  <= 20'h42442; 
			12'd1252 :q  <= 20'h7b824; 
			12'd1253 :q  <= 20'h1b042; 
			12'd1254 :q  <= 20'h63c42; 
			12'd1255 :q  <= 20'h4b442; 
			12'd1256 :q  <= 20'h22dc9; 
			12'd1257 :q  <= 20'h3b483; 
			12'd1258 :q  <= 20'h7b824; 
			12'd1259 :q  <= 20'h23824; 
			12'd1260 :q  <= 20'h700cd; 
			12'd1261 :q  <= 20'h2044c; 
			12'd1262 :q  <= 20'h5b8c6; 
			12'd1263 :q  <= 20'h1b8c6; 
			12'd1264 :q  <= 20'h74462; 
			12'd1265 :q  <= 20'h1c462; 
			12'd1266 :q  <= 20'h700cd; 
			12'd1267 :q  <= 20'h000cd; 
			12'd1268 :q  <= 20'h528e6; 
			12'd1269 :q  <= 20'h33c42; 
			12'd1270 :q  <= 20'h32d06; 
			12'd1271 :q  <= 20'h39842; 
			12'd1272 :q  <= 20'h10a06; 
			12'd1273 :q  <= 20'h29063; 
			12'd1274 :q  <= 20'h59c6a; 
			12'd1275 :q  <= 20'h31c6a; 
			12'd1276 :q  <= 20'h51c62; 
			12'd1277 :q  <= 20'h43082; 
			12'd1278 :q  <= 20'h50423; 
			12'd1279 :q  <= 20'h08892; 
			12'd1280 :q  <= 20'h6108c; 
			12'd1281 :q  <= 20'h00026; 
			12'd1282 :q  <= 20'h4ac43; 
			12'd1283 :q  <= 20'h41c83; 
			12'd1284 :q  <= 20'h51c62; 
			12'd1285 :q  <= 20'h39c62; 
			12'd1286 :q  <= 20'h490c1; 
			12'd1287 :q  <= 20'h41c43; 
			12'd1288 :q  <= 20'h61d06; 
			12'd1289 :q  <= 20'h01d06; 
			12'd1290 :q  <= 20'h9084a; 
			12'd1291 :q  <= 20'h008c4; 
			12'd1292 :q  <= 20'h490c1; 
			12'd1293 :q  <= 20'h3bc42; 
			12'd1294 :q  <= 20'h5b426; 
			12'd1295 :q  <= 20'h43426; 
			12'd1296 :q  <= 20'h70c41; 
			12'd1297 :q  <= 20'h43c43; 
			12'd1298 :q  <= 20'h63ce4; 
			12'd1299 :q  <= 20'h23983; 
			12'd1300 :q  <= 20'h50c62; 
			12'd1301 :q  <= 20'h23042; 
			12'd1302 :q  <= 20'h52c86; 
			12'd1303 :q  <= 20'h3b442; 
			12'd1304 :q  <= 20'h22dc4; 
			12'd1305 :q  <= 20'h0ca42; 
			12'd1306 :q  <= 20'h5c842; 
			12'd1307 :q  <= 20'h3c842; 
			12'd1308 :q  <= 20'h64902; 
			12'd1309 :q  <= 20'h3b8c2; 
			12'd1310 :q  <= 20'h43088; 
			12'd1311 :q  <= 20'h22463; 
			12'd1312 :q  <= 20'h3a8c2; 
			12'd1313 :q  <= 20'h2808f; 
			12'd1314 :q  <= 20'h4198e; 
			12'd1315 :q  <= 20'h2c063; 
			12'd1316 :q  <= 20'h40593; 
			12'd1317 :q  <= 20'h18062; 
			12'd1318 :q  <= 20'h53085; 
			12'd1319 :q  <= 20'h33085; 
			12'd1320 :q  <= 20'h5ac42; 
			12'd1321 :q  <= 20'h00866; 
			12'd1322 :q  <= 20'h5ac42; 
			12'd1323 :q  <= 20'h3988a; 
			12'd1324 :q  <= 20'h5ac42; 
			12'd1325 :q  <= 20'h134a2; 
			12'd1326 :q  <= 20'h5ac42; 
			12'd1327 :q  <= 20'h3ac42; 
			12'd1328 :q  <= 20'h73463; 
			12'd1329 :q  <= 20'h1b463; 
			12'd1330 :q  <= 20'h4b843; 
			12'd1331 :q  <= 20'h41c63; 
			12'd1332 :q  <= 20'h69463; 
			12'd1333 :q  <= 20'h024a3; 
			12'd1334 :q  <= 20'h69463; 
			12'd1335 :q  <= 20'h4b048; 
			12'd1336 :q  <= 20'h59c42; 
			12'd1337 :q  <= 20'h040c4; 
			12'd1338 :q  <= 20'h51843; 
			12'd1339 :q  <= 20'h49446; 
			12'd1340 :q  <= 20'h63d04; 
			12'd1341 :q  <= 20'h03906; 
			12'd1342 :q  <= 20'h48062; 
			12'd1343 :q  <= 20'h23c82; 
			12'd1344 :q  <= 20'h61c6d; 
			12'd1345 :q  <= 20'h29c6d; 
			12'd1346 :q  <= 20'h49869; 
			12'd1347 :q  <= 20'h210ec; 
			12'd1348 :q  <= 20'h63042; 
			12'd1349 :q  <= 20'h33042; 
			12'd1350 :q  <= 20'h42482; 
			12'd1351 :q  <= 20'h19842; 
			12'd1352 :q  <= 20'h81862; 
			12'd1353 :q  <= 20'h01e64; 
			12'd1354 :q  <= 20'h50941; 
			12'd1355 :q  <= 20'h4904c; 
			12'd1356 :q  <= 20'h64881; 
			12'd1357 :q  <= 20'h09cc4; 
			12'd1358 :q  <= 20'h600cd; 
			12'd1359 :q  <= 20'h100cd; 
			12'd1360 :q  <= 20'h51508; 
			12'd1361 :q  <= 20'h40c45; 
			12'd1362 :q  <= 20'h41121; 
			12'd1363 :q  <= 20'h19121; 
			12'd1364 :q  <= 20'h0824a; 
			12'd1365 :q  <= 20'h3c4a3; 
			12'd1366 :q  <= 20'h3acc1; 
			12'd1367 :q  <= 20'h10862; 
			12'd1368 :q  <= 20'h43082; 
			12'd1369 :q  <= 20'h32866; 
			12'd1370 :q  <= 20'h59044; 
			12'd1371 :q  <= 20'h39044; 
			12'd1372 :q  <= 20'h49844; 
			12'd1373 :q  <= 20'h33503; 
			12'd1374 :q  <= 20'h4bc64; 
			12'd1375 :q  <= 20'h48851; 
			12'd1376 :q  <= 20'h380c1; 
			12'd1377 :q  <= 20'h43c64; 
			12'd1378 :q  <= 20'h3b4e3; 
			12'd1379 :q  <= 20'h44063; 
			12'd1380 :q  <= 20'h3090a; 
			12'd1381 :q  <= 20'h11508; 
			12'd1382 :q  <= 20'h74042; 
			12'd1383 :q  <= 20'h24042; 
			12'd1384 :q  <= 20'h52c86; 
			12'd1385 :q  <= 20'h32c86; 
			12'd1386 :q  <= 20'h53823; 
			12'd1387 :q  <= 20'h43883; 
			12'd1388 :q  <= 20'h50086; 
			12'd1389 :q  <= 20'h00e82; 
			12'd1390 :q  <= 20'h60102; 
			12'd1391 :q  <= 20'h13148; 
			12'd1392 :q  <= 20'h89c4a; 
			12'd1393 :q  <= 20'h09c4a; 
			12'd1394 :q  <= 20'h7a866; 
			12'd1395 :q  <= 20'h210c2; 
			12'd1396 :q  <= 20'h01686; 
			12'd1397 :q  <= 20'h00102; 
			12'd1398 :q  <= 20'h08244; 
			12'd1399 :q  <= 20'h0b4c2; 
			12'd1400 :q  <= 20'h52064; 
			12'd1401 :q  <= 20'h304c1; 
			12'd1402 :q  <= 20'h43883; 
			12'd1403 :q  <= 20'h09a42; 
			12'd1404 :q  <= 20'h7ac22; 
			12'd1405 :q  <= 20'h31422; 
			12'd1406 :q  <= 20'h69023; 
			12'd1407 :q  <= 20'h13c22; 
			12'd1408 :q  <= 20'h61083; 
			12'd1409 :q  <= 20'h000e3; 
			12'd1410 :q  <= 20'h4b0c2; 
			12'd1411 :q  <= 20'h29043; 
			12'd1412 :q  <= 20'h91043; 
			12'd1413 :q  <= 20'h18106; 
			12'd1414 :q  <= 20'h00a86; 
			12'd1415 :q  <= 20'h21c44; 
			12'd1416 :q  <= 20'h1a9e2; 
			12'd1417 :q  <= 20'h1818b; 
			12'd1418 :q  <= 20'h68046; 
			12'd1419 :q  <= 20'h04c41; 
			12'd1420 :q  <= 20'h8288a; 
			12'd1421 :q  <= 20'h22143; 
			12'd1422 :q  <= 20'h73063; 
			12'd1423 :q  <= 20'h0288a; 
			12'd1424 :q  <= 20'h90c46; 
			12'd1425 :q  <= 20'h31823; 
			12'd1426 :q  <= 20'h39ce2; 
			12'd1427 :q  <= 20'h00c46; 
			12'd1428 :q  <= 20'h58461; 
			12'd1429 :q  <= 20'h28046; 
			12'd1430 :q  <= 20'h0864e; 
			12'd1431 :q  <= 20'h21903; 
			12'd1432 :q  <= 20'h4b0c2; 
			12'd1433 :q  <= 20'h2b0c2; 
			12'd1434 :q  <= 20'h51c65; 
			12'd1435 :q  <= 20'h39c65; 
			12'd1436 :q  <= 20'h6806a; 
			12'd1437 :q  <= 20'h22c62; 
			12'd1438 :q  <= 20'h88c66; 
			12'd1439 :q  <= 20'h0a24a; 
			12'd1440 :q  <= 20'h6806a; 
			12'd1441 :q  <= 20'h4b843; 
			12'd1442 :q  <= 20'h80c67; 
			12'd1443 :q  <= 20'h2006a; 
			12'd1444 :q  <= 20'h80c67; 
			12'd1445 :q  <= 20'h02422; 
			12'd1446 :q  <= 20'h9044a; 
			12'd1447 :q  <= 20'h0044a; 
			12'd1448 :q  <= 20'h54064; 
			12'd1449 :q  <= 20'h12063; 
			12'd1450 :q  <= 20'h58046; 
			12'd1451 :q  <= 20'h38046; 
			12'd1452 :q  <= 20'h80c67; 
			12'd1453 :q  <= 20'h08c67; 
			12'd1454 :q  <= 20'h704d0; 
			12'd1455 :q  <= 20'h004d0; 
			12'd1456 :q  <= 20'h10208; 
			12'd1457 :q  <= 20'h320a3; 
			12'd1458 :q  <= 20'h49c63; 
			12'd1459 :q  <= 20'h42083; 
			12'd1460 :q  <= 20'h49844; 
			12'd1461 :q  <= 20'h01de1; 
			12'd1462 :q  <= 20'h408e9; 
			12'd1463 :q  <= 20'h09e04; 
			12'd1464 :q  <= 20'h33102; 
			12'd1465 :q  <= 20'h42c63; 
			12'd1466 :q  <= 20'h215ca; 
			12'd1467 :q  <= 20'h23062; 
			12'd1468 :q  <= 20'h4acc1; 
			12'd1469 :q  <= 20'h224e6; 
			12'd1470 :q  <= 20'h3a8c3; 
			12'd1471 :q  <= 20'h4ac42; 
			12'd1472 :q  <= 20'h01686; 
			12'd1473 :q  <= 20'h310c1; 
			12'd1474 :q  <= 20'h4acc1; 
			12'd1475 :q  <= 20'h2acc1; 
			12'd1476 :q  <= 20'h54064; 
			12'd1477 :q  <= 20'h41c63; 
			12'd1478 :q  <= 20'h13208; 
			12'd1479 :q  <= 20'h03de2; 
			12'd1480 :q  <= 20'h790a6; 
			12'd1481 :q  <= 20'h49444; 
			12'd1482 :q  <= 20'h42926; 
			12'd1483 :q  <= 20'h14de1; 
			12'd1484 :q  <= 20'h54064; 
			12'd1485 :q  <= 20'h03e84; 
			12'd1486 :q  <= 20'h54064; 
			12'd1487 :q  <= 20'h3c064; 
			12'd1488 :q  <= 20'h4c063; 
			12'd1489 :q  <= 20'h42c86; 
			12'd1490 :q  <= 20'h4984c; 
			12'd1491 :q  <= 20'h44483; 
			12'd1492 :q  <= 20'h4c902; 
			12'd1493 :q  <= 20'h0c902; 
			12'd1494 :q  <= 20'h694cf; 
			12'd1495 :q  <= 20'h4a042; 
			12'd1496 :q  <= 20'h49443; 
			12'd1497 :q  <= 20'h094cf; 
			12'd1498 :q  <= 20'h205c8; 
			12'd1499 :q  <= 20'h11090; 
			12'd1500 :q  <= 20'h6106c; 
			12'd1501 :q  <= 20'h2154c; 
			12'd1502 :q  <= 20'h4b843; 
			12'd1503 :q  <= 20'h29043; 
			12'd1504 :q  <= 20'h6088a; 
			12'd1505 :q  <= 20'h310e3; 
			12'd1506 :q  <= 20'h10242; 
			12'd1507 :q  <= 20'h00242; 
			12'd1508 :q  <= 20'h6b486; 
			12'd1509 :q  <= 20'h1b486; 
			12'd1510 :q  <= 20'h53046; 
			12'd1511 :q  <= 20'h2a54a; 
			12'd1512 :q  <= 20'h59082; 
			12'd1513 :q  <= 20'h3b0c8; 
			12'd1514 :q  <= 20'h6088a; 
			12'd1515 :q  <= 20'h42c41; 
			12'd1516 :q  <= 20'h5142c; 
			12'd1517 :q  <= 20'h02cc9; 
			12'd1518 :q  <= 20'h6088a; 
			12'd1519 :q  <= 20'h2088a; 
			12'd1520 :q  <= 20'h59082; 
			12'd1521 :q  <= 20'h038c3; 
			12'd1522 :q  <= 20'h59082; 
			12'd1523 :q  <= 20'h30462; 
			12'd1524 :q  <= 20'h59082; 
			12'd1525 :q  <= 20'h29082; 
			12'd1526 :q  <= 20'h6804c; 
			12'd1527 :q  <= 20'h3006a; 
			12'd1528 :q  <= 20'h18228; 
			12'd1529 :q  <= 20'h01284; 
			12'd1530 :q  <= 20'h00d02; 
			12'd1531 :q  <= 20'h42c83; 
			12'd1532 :q  <= 20'h29cc4; 
			12'd1533 :q  <= 20'h40c89; 
			12'd1534 :q  <= 20'h43c24; 
			12'd1535 :q  <= 20'h21587; 
			12'd1536 :q  <= 20'h2088a; 
			12'd1537 :q  <= 20'h18222; 
			12'd1538 :q  <= 20'h10a0f; 
			12'd1539 :q  <= 20'h788a2; 
			12'd1540 :q  <= 20'h48c42; 
			12'd1541 :q  <= 20'h2160f; 
			12'd1542 :q  <= 20'h3b4a6; 
			12'd1543 :q  <= 20'h51c62; 
			12'd1544 :q  <= 20'h40c61; 
			12'd1545 :q  <= 20'h4c063; 
			12'd1546 :q  <= 20'h008a2; 
			12'd1547 :q  <= 20'h61483; 
			12'd1548 :q  <= 20'h09d81; 
			12'd1549 :q  <= 20'h394ce; 
			12'd1550 :q  <= 20'h0010a; 
			12'd1551 :q  <= 20'h48462; 
			12'd1552 :q  <= 20'h40462; 
			12'd1553 :q  <= 20'h61063; 
			12'd1554 :q  <= 20'h390d0; 
			12'd1555 :q  <= 20'h61063; 
			12'd1556 :q  <= 20'h10c46; 
			12'd1557 :q  <= 20'h708c9; 
			12'd1558 :q  <= 20'h29063; 
			12'd1559 :q  <= 20'h4c462; 
			12'd1560 :q  <= 20'h29443; 
			12'd1561 :q  <= 20'h6ac66; 
			12'd1562 :q  <= 20'h1b846; 
			12'd1563 :q  <= 20'h70cc2; 
			12'd1564 :q  <= 20'h02202; 
			12'd1565 :q  <= 20'h70cc2; 
			12'd1566 :q  <= 20'h000a6; 
			12'd1567 :q  <= 20'h61483; 
			12'd1568 :q  <= 20'h22c66; 
			12'd1569 :q  <= 20'h61483; 
			12'd1570 :q  <= 20'h49423; 
			12'd1571 :q  <= 20'h61483; 
			12'd1572 :q  <= 20'h3190c; 
			12'd1573 :q  <= 20'h61483; 
			12'd1574 :q  <= 20'h2b122; 
			12'd1575 :q  <= 20'h61483; 
			12'd1576 :q  <= 20'h21483; 
			12'd1577 :q  <= 20'h31922; 
			12'd1578 :q  <= 20'h22c23; 
			12'd1579 :q  <= 20'h730c6; 
			12'd1580 :q  <= 20'h38067; 
			12'd1581 :q  <= 20'h4a063; 
			12'd1582 :q  <= 20'h42063; 
			12'd1583 :q  <= 20'h2a963; 
			12'd1584 :q  <= 20'h29d41; 
			12'd1585 :q  <= 20'h49c62; 
			12'd1586 :q  <= 20'h41c62; 
			12'd1587 :q  <= 20'h5a482; 
			12'd1588 :q  <= 20'h2a482; 
			12'd1589 :q  <= 20'h72844; 
			12'd1590 :q  <= 20'h39c62; 
			12'd1591 :q  <= 20'h744c3; 
			12'd1592 :q  <= 20'h2158c; 
			12'd1593 :q  <= 20'h32508; 
			12'd1594 :q  <= 20'h011e4; 
			12'd1595 :q  <= 20'h68881; 
			12'd1596 :q  <= 20'h23042; 
			12'd1597 :q  <= 20'h43483; 
			12'd1598 :q  <= 20'h4b443; 
			12'd1599 :q  <= 20'h6ac43; 
			12'd1600 :q  <= 20'h3b084; 
			12'd1601 :q  <= 20'h52c42; 
			12'd1602 :q  <= 20'h44462; 
			12'd1603 :q  <= 20'h52c42; 
			12'd1604 :q  <= 20'h044c3; 
			12'd1605 :q  <= 20'h52c42; 
			12'd1606 :q  <= 20'h42c42; 
			12'd1607 :q  <= 20'h61504; 
			12'd1608 :q  <= 20'h01504; 
			12'd1609 :q  <= 20'h68881; 
			12'd1610 :q  <= 20'h18881; 
			12'd1611 :q  <= 20'h50082; 
			12'd1612 :q  <= 20'h3b061; 
			12'd1613 :q  <= 20'h42c88; 
			12'd1614 :q  <= 20'h4a442; 
			12'd1615 :q  <= 20'h1c9e2; 
			12'd1616 :q  <= 20'h1184c; 
			12'd1617 :q  <= 20'h4a043; 
			12'd1618 :q  <= 20'h3a862; 
			12'd1619 :q  <= 20'h5ac61; 
			12'd1620 :q  <= 20'h32c61; 
			12'd1621 :q  <= 20'h48882; 
			12'd1622 :q  <= 20'h23043; 
			12'd1623 :q  <= 20'h10643; 
			12'd1624 :q  <= 20'h2848e; 
			12'd1625 :q  <= 20'h44183; 
			12'd1626 :q  <= 20'h0c643; 
			12'd1627 :q  <= 20'h4b846; 
			12'd1628 :q  <= 20'h4b028; 
			12'd1629 :q  <= 20'h4b843; 
			12'd1630 :q  <= 20'h4984c; 
			12'd1631 :q  <= 20'h62463; 
			12'd1632 :q  <= 20'h00488; 
			12'd1633 :q  <= 20'h484c2; 
			12'd1634 :q  <= 20'h08d8e; 
			12'd1635 :q  <= 20'h43082; 
			12'd1636 :q  <= 20'h0a542; 
			12'd1637 :q  <= 20'h43c83; 
			12'd1638 :q  <= 20'h32103; 
			12'd1639 :q  <= 20'h4bca3; 
			12'd1640 :q  <= 20'h41c83; 
			12'd1641 :q  <= 20'h39cc2; 
			12'd1642 :q  <= 20'h29d02; 
			12'd1643 :q  <= 20'h62463; 
			12'd1644 :q  <= 20'h21c82; 
			12'd1645 :q  <= 20'h708c9; 
			12'd1646 :q  <= 20'h22463; 
			12'd1647 :q  <= 20'h62463; 
			12'd1648 :q  <= 20'h008c9; 
			12'd1649 :q  <= 20'h88c66; 
			12'd1650 :q  <= 20'h00c66; 
			12'd1651 :q  <= 20'h8b822; 
			12'd1652 :q  <= 20'h22483; 
			12'd1653 :q  <= 20'h62463; 
			12'd1654 :q  <= 20'h2a463; 
			12'd1655 :q  <= 20'h494c8; 
			12'd1656 :q  <= 20'h294c8; 
			12'd1657 :q  <= 20'h80486; 
			12'd1658 :q  <= 20'h080d4; 
			12'd1659 :q  <= 20'h62c62; 
			12'd1660 :q  <= 20'h2ac62; 
			12'd1661 :q  <= 20'h490c1; 
			12'd1662 :q  <= 20'h00103; 
			12'd1663 :q  <= 20'h78045; 
			12'd1664 :q  <= 20'h20462; 
			12'd1665 :q  <= 20'h380cf; 
			12'd1666 :q  <= 20'h32c61; 
			12'd1667 :q  <= 20'h60064; 
			12'd1668 :q  <= 20'h290c1; 
			12'd1669 :q  <= 20'h61c62; 
			12'd1670 :q  <= 20'h00486; 
			12'd1671 :q  <= 20'h61c62; 
			12'd1672 :q  <= 20'h14063; 
			12'd1673 :q  <= 20'h6a0ca; 
			12'd1674 :q  <= 20'h024a2; 
			12'd1675 :q  <= 20'h62c42; 
			12'd1676 :q  <= 20'h1bc63; 
			12'd1677 :q  <= 20'h61c62; 
			12'd1678 :q  <= 20'h29c62; 
			12'd1679 :q  <= 20'h49529; 
			12'd1680 :q  <= 20'h28067; 
			12'd1681 :q  <= 20'h28985; 
			12'd1682 :q  <= 20'h32c42; 
			12'd1683 :q  <= 20'h7bc62; 
			12'd1684 :q  <= 20'h13c62; 
			12'd1685 :q  <= 20'h730c8; 
			12'd1686 :q  <= 20'h121e6; 
			12'd1687 :q  <= 20'h10a51; 
			12'd1688 :q  <= 20'h28481; 
			12'd1689 :q  <= 20'h28985; 
			12'd1690 :q  <= 20'h18985; 
			12'd1691 :q  <= 20'h22584; 
			12'd1692 :q  <= 20'h2bcc2; 
			12'd1693 :q  <= 20'h53843; 
			12'd1694 :q  <= 20'h03682; 
			12'd1695 :q  <= 20'h22588; 
			12'd1696 :q  <= 20'h43466; 
			12'd1697 :q  <= 20'h53042; 
			12'd1698 :q  <= 20'h4b042; 
			12'd1699 :q  <= 20'h22dc4; 
			12'd1700 :q  <= 20'h41482; 
			12'd1701 :q  <= 20'h528c3; 
			12'd1702 :q  <= 20'h13822; 
			12'd1703 :q  <= 20'h6a0cc; 
			12'd1704 :q  <= 20'h0a0cc; 
			12'd1705 :q  <= 20'h500ca; 
			12'd1706 :q  <= 20'h2ad04; 
			12'd1707 :q  <= 20'h54104; 
			12'd1708 :q  <= 20'h39cc6; 
			12'd1709 :q  <= 20'h5088a; 
			12'd1710 :q  <= 20'h30489; 
			12'd1711 :q  <= 20'h64c41; 
			12'd1712 :q  <= 20'h08889; 
			12'd1713 :q  <= 20'h394c4; 
			12'd1714 :q  <= 20'h49044; 
			12'd1715 :q  <= 20'h71448; 
			12'd1716 :q  <= 20'h398ac; 
			12'd1717 :q  <= 20'h71846; 
			12'd1718 :q  <= 20'h21846; 
			12'd1719 :q  <= 20'h43d44; 
			12'd1720 :q  <= 20'h34842; 
			12'd1721 :q  <= 20'h58cc2; 
			12'd1722 :q  <= 20'h10206; 
			12'd1723 :q  <= 20'h58cc2; 
			12'd1724 :q  <= 20'h22d43; 
			12'd1725 :q  <= 20'h58cc2; 
			12'd1726 :q  <= 20'h18cc2; 
			12'd1727 :q  <= 20'h80087; 
			12'd1728 :q  <= 20'h03926; 
			12'd1729 :q  <= 20'h4c063; 
			12'd1730 :q  <= 20'h218c2; 
			12'd1731 :q  <= 20'h7ac23; 
			12'd1732 :q  <= 20'h29443; 
			12'd1733 :q  <= 20'h52442; 
			12'd1734 :q  <= 20'h18483; 
			12'd1735 :q  <= 20'h80087; 
			12'd1736 :q  <= 20'h00281; 
			12'd1737 :q  <= 20'h7ac23; 
			12'd1738 :q  <= 20'h01064; 
			12'd1739 :q  <= 20'h80c66; 
			12'd1740 :q  <= 20'h08c66; 
			12'd1741 :q  <= 20'h30986; 
			12'd1742 :q  <= 20'h42883; 
			12'd1743 :q  <= 20'h209c6; 
			12'd1744 :q  <= 20'h4ac43; 
			12'd1745 :q  <= 20'h7b443; 
			12'd1746 :q  <= 20'h43083; 
			12'd1747 :q  <= 20'h7ac23; 
			12'd1748 :q  <= 20'h3b4a2; 
			12'd1749 :q  <= 20'h3b0c3; 
			12'd1750 :q  <= 20'h2ac84; 
			12'd1751 :q  <= 20'h59063; 
			12'd1752 :q  <= 20'h31063; 
			12'd1753 :q  <= 20'h81466; 
			12'd1754 :q  <= 20'h19987; 
			12'd1755 :q  <= 20'h81466; 
			12'd1756 :q  <= 20'h1b443; 
			12'd1757 :q  <= 20'h81466; 
			12'd1758 :q  <= 20'h09466; 
			12'd1759 :q  <= 20'h0a641; 
			12'd1760 :q  <= 20'h02507; 
			12'd1761 :q  <= 20'h62d02; 
			12'd1762 :q  <= 20'h02d02; 
			12'd1763 :q  <= 20'h4b443; 
			12'd1764 :q  <= 20'h22984; 
			12'd1765 :q  <= 20'h48c67; 
			12'd1766 :q  <= 20'h38865; 
			12'd1767 :q  <= 20'h4b086; 
			12'd1768 :q  <= 20'h41c66; 
			12'd1769 :q  <= 20'h79082; 
			12'd1770 :q  <= 20'h41c63; 
			12'd1771 :q  <= 20'h708c4; 
			12'd1772 :q  <= 20'h3c0c1; 
			12'd1773 :q  <= 20'h7b443; 
			12'd1774 :q  <= 20'h41c6a; 
			12'd1775 :q  <= 20'h5a846; 
			12'd1776 :q  <= 20'h32881; 
			12'd1777 :q  <= 20'h52442; 
			12'd1778 :q  <= 20'h42442; 
			12'd1779 :q  <= 20'h61c42; 
			12'd1780 :q  <= 20'h29c42; 
			12'd1781 :q  <= 20'h6806e; 
			12'd1782 :q  <= 20'h2006e; 
			12'd1783 :q  <= 20'h6906e; 
			12'd1784 :q  <= 20'h4b843; 
			12'd1785 :q  <= 20'h43883; 
			12'd1786 :q  <= 20'h20870; 
			12'd1787 :q  <= 20'h3890a; 
			12'd1788 :q  <= 20'h338e3; 
			12'd1789 :q  <= 20'h4894c; 
			12'd1790 :q  <= 20'h31d02; 
			12'd1791 :q  <= 20'h43486; 
			12'd1792 :q  <= 20'h31823; 
			12'd1793 :q  <= 20'h80886; 
			12'd1794 :q  <= 20'h31882; 
			12'd1795 :q  <= 20'h80886; 
			12'd1796 :q  <= 20'h00886; 
			12'd1797 :q  <= 20'h49846; 
			12'd1798 :q  <= 20'h190ca; 
			12'd1799 :q  <= 20'h49446; 
			12'd1800 :q  <= 20'h1b443; 
			12'd1801 :q  <= 20'h6b462; 
			12'd1802 :q  <= 20'h14144; 
			12'd1803 :q  <= 20'h29946; 
			12'd1804 :q  <= 20'h3b823; 
			12'd1805 :q  <= 20'h740c3; 
			12'd1806 :q  <= 20'h29063; 
			12'd1807 :q  <= 20'h39143; 
			12'd1808 :q  <= 20'h010a4; 
			12'd1809 :q  <= 20'h6ac69; 
			12'd1810 :q  <= 20'h22c69; 
			12'd1811 :q  <= 20'h49c41; 
			12'd1812 :q  <= 20'h280d1; 
			12'd1813 :q  <= 20'h50cc3; 
			12'd1814 :q  <= 20'h109e4; 
			12'd1815 :q  <= 20'h40902; 
			12'd1816 :q  <= 20'h40466; 
			12'd1817 :q  <= 20'h4c442; 
			12'd1818 :q  <= 20'h0004e; 
			12'd1819 :q  <= 20'h600e3; 
			12'd1820 :q  <= 20'h0b822; 
			12'd1821 :q  <= 20'h73048; 
			12'd1822 :q  <= 20'h080e3; 
			12'd1823 :q  <= 20'h73048; 
			12'd1824 :q  <= 20'h3010c; 
			12'd1825 :q  <= 20'h30509; 
			12'd1826 :q  <= 20'h28842; 
			12'd1827 :q  <= 20'h6b8c6; 
			12'd1828 :q  <= 20'h04682; 
			12'd1829 :q  <= 20'h50c46; 
			12'd1830 :q  <= 20'h2b0c2; 
			12'd1831 :q  <= 20'h51ccd; 
			12'd1832 :q  <= 20'h2bd45; 
			12'd1833 :q  <= 20'h5108a; 
			12'd1834 :q  <= 20'h29c41; 
			12'd1835 :q  <= 20'h50cc7; 
			12'd1836 :q  <= 20'h20cc7; 
			12'd1837 :q  <= 20'h09e45; 
			12'd1838 :q  <= 20'h1c483; 
			12'd1839 :q  <= 20'h43986; 
			12'd1840 :q  <= 20'h03684; 
			12'd1841 :q  <= 20'h215c2; 
			12'd1842 :q  <= 20'h0894c; 
			12'd1843 :q  <= 20'h305c3; 
			12'd1844 :q  <= 20'h44043; 
			12'd1845 :q  <= 20'h4c462; 
			12'd1846 :q  <= 20'h2bc82; 
			12'd1847 :q  <= 20'h53c23; 
			12'd1848 :q  <= 20'h44084; 
			12'd1849 :q  <= 20'h32d06; 
			12'd1850 :q  <= 20'h134a2; 
			12'd1851 :q  <= 20'h6b8c6; 
			12'd1852 :q  <= 20'h0a644; 
			12'd1853 :q  <= 20'h6b8c6; 
			12'd1854 :q  <= 20'h00826; 
			12'd1855 :q  <= 20'h281f4; 
			12'd1856 :q  <= 20'h0b8c6; 
			12'd1857 :q  <= 20'h43886; 
			12'd1858 :q  <= 20'h3ac41; 
			12'd1859 :q  <= 20'h4c462; 
			12'd1860 :q  <= 20'h44462; 
			12'd1861 :q  <= 20'h63886; 
			12'd1862 :q  <= 20'h23886; 
			12'd1863 :q  <= 20'h6b846; 
			12'd1864 :q  <= 20'h2b846; 
			12'd1865 :q  <= 20'h380cc; 
			12'd1866 :q  <= 20'h01d82; 
			12'd1867 :q  <= 20'h50c6d; 
			12'd1868 :q  <= 20'h38c6d; 
			12'd1869 :q  <= 20'h520c3; 
			12'd1870 :q  <= 20'h1ac62; 
			12'd1871 :q  <= 20'h6b0c8; 
			12'd1872 :q  <= 20'h398c5; 
			12'd1873 :q  <= 20'h8ac47; 
			12'd1874 :q  <= 20'h1b502; 
			12'd1875 :q  <= 20'h32503; 
			12'd1876 :q  <= 20'h20c83; 
			12'd1877 :q  <= 20'h58c83; 
			12'd1878 :q  <= 20'h0922c; 
			12'd1879 :q  <= 20'h58c83; 
			12'd1880 :q  <= 20'h220c3; 
			12'd1881 :q  <= 20'h60ca3; 
			12'd1882 :q  <= 20'h0ac47; 
			12'd1883 :q  <= 20'h7b048; 
			12'd1884 :q  <= 20'h22163; 
			12'd1885 :q  <= 20'h4b4c2; 
			12'd1886 :q  <= 20'h33483; 
			12'd1887 :q  <= 20'h4b063; 
			12'd1888 :q  <= 20'h28c63; 
			12'd1889 :q  <= 20'h49043; 
			12'd1890 :q  <= 20'h00a03; 
			12'd1891 :q  <= 20'h7b048; 
			12'd1892 :q  <= 20'h1b048; 
			12'd1893 :q  <= 20'h73466; 
			12'd1894 :q  <= 20'h1b466; 
			12'd1895 :q  <= 20'h31542; 
			12'd1896 :q  <= 20'h139c6; 
			12'd1897 :q  <= 20'h53823; 
			12'd1898 :q  <= 20'h24042; 
			12'd1899 :q  <= 20'h51843; 
			12'd1900 :q  <= 20'h04682; 
			12'd1901 :q  <= 20'h69823; 
			12'd1902 :q  <= 20'h43462; 
			12'd1903 :q  <= 20'h60863; 
			12'd1904 :q  <= 20'h1c842; 
			12'd1905 :q  <= 20'h4c064; 
			12'd1906 :q  <= 20'h31823; 
			12'd1907 :q  <= 20'h684a2; 
			12'd1908 :q  <= 20'h3b8c2; 
			12'd1909 :q  <= 20'h58c64; 
			12'd1910 :q  <= 20'h0b586; 
			12'd1911 :q  <= 20'h72ca2; 
			12'd1912 :q  <= 20'h13dc4; 
			12'd1913 :q  <= 20'h19dc2; 
			12'd1914 :q  <= 20'h0ac82; 
			12'd1915 :q  <= 20'h700ce; 
			12'd1916 :q  <= 20'h22c23; 
			12'd1917 :q  <= 20'h700ce; 
			12'd1918 :q  <= 20'h0a867; 
			12'd1919 :q  <= 20'h43122; 
			12'd1920 :q  <= 20'h01a81; 
			12'd1921 :q  <= 20'h41084; 
			12'd1922 :q  <= 20'h00042; 
			12'd1923 :q  <= 20'h28d49; 
			12'd1924 :q  <= 20'h7888a; 
			12'd1925 :q  <= 20'h40847; 
			12'd1926 :q  <= 20'h39181; 
			12'd1927 :q  <= 20'h19121; 
			12'd1928 :q  <= 20'h7a824; 
			12'd1929 :q  <= 20'h228c4; 
			12'd1930 :q  <= 20'h7a426; 
			12'd1931 :q  <= 20'h3c4c3; 
			12'd1932 :q  <= 20'h70c50; 
			12'd1933 :q  <= 20'h22426; 
			12'd1934 :q  <= 20'h604a2; 
			12'd1935 :q  <= 20'h34882; 
			12'd1936 :q  <= 20'h1120a; 
			12'd1937 :q  <= 20'h3142a; 
			12'd1938 :q  <= 20'h221e2; 
			12'd1939 :q  <= 20'h0a1e2; 
			12'd1940 :q  <= 20'h49466; 
			12'd1941 :q  <= 20'h29d02; 
			12'd1942 :q  <= 20'h4ac43; 
			12'd1943 :q  <= 20'h08203; 
			12'd1944 :q  <= 20'h588e2; 
			12'd1945 :q  <= 20'h28552; 
			12'd1946 :q  <= 20'h89062; 
			12'd1947 :q  <= 20'h43423; 
			12'd1948 :q  <= 20'h1b9c6; 
			12'd1949 :q  <= 20'h00864; 
			12'd1950 :q  <= 20'h604a2; 
			12'd1951 :q  <= 20'h184a2; 
			12'd1952 :q  <= 20'h53443; 
			12'd1953 :q  <= 20'h43443; 
			12'd1954 :q  <= 20'h73043; 
			12'd1955 :q  <= 20'h38843; 
			12'd1956 :q  <= 20'h29944; 
			12'd1957 :q  <= 20'h4b426; 
			12'd1958 :q  <= 20'h53042; 
			12'd1959 :q  <= 20'h23043; 
			12'd1960 :q  <= 20'h710c6; 
			12'd1961 :q  <= 20'h44443; 
			12'd1962 :q  <= 20'h81086; 
			12'd1963 :q  <= 20'h01086; 
			12'd1964 :q  <= 20'h71843; 
			12'd1965 :q  <= 20'h22501; 
			12'd1966 :q  <= 20'h43083; 
			12'd1967 :q  <= 20'h2b146; 
			12'd1968 :q  <= 20'h5b022; 
			12'd1969 :q  <= 20'h43c82; 
			12'd1970 :q  <= 20'h32508; 
			12'd1971 :q  <= 20'h3b086; 
			12'd1972 :q  <= 20'h52c61; 
			12'd1973 :q  <= 20'h49c4a; 
			12'd1974 :q  <= 20'h400c6; 
			12'd1975 :q  <= 20'h1ac46; 
			12'd1976 :q  <= 20'h83022; 
			12'd1977 :q  <= 20'h0b8c6; 
			12'd1978 :q  <= 20'h68466; 
			12'd1979 :q  <= 20'h42042; 
			12'd1980 :q  <= 20'h4a463; 
			12'd1981 :q  <= 20'h41c63; 
			12'd1982 :q  <= 20'h70043; 
			12'd1983 :q  <= 20'h08249; 
			12'd1984 :q  <= 20'h5948f; 
			12'd1985 :q  <= 20'h2948f; 
			12'd1986 :q  <= 20'h70043; 
			12'd1987 :q  <= 20'h20043; 
			12'd1988 :q  <= 20'h5b042; 
			12'd1989 :q  <= 20'h3b042; 
			12'd1990 :q  <= 20'h60064; 
			12'd1991 :q  <= 20'h22c63; 
			12'd1992 :q  <= 20'h61c82; 
			12'd1993 :q  <= 20'h42862; 
			12'd1994 :q  <= 20'h4a462; 
			12'd1995 :q  <= 20'h42462; 
			12'd1996 :q  <= 20'h60064; 
			12'd1997 :q  <= 20'h28064; 
			12'd1998 :q  <= 20'h23984; 
			12'd1999 :q  <= 20'h43443; 
			12'd2000 :q  <= 20'h52868; 
			12'd2001 :q  <= 20'h42888; 
			12'd2002 :q  <= 20'h52061; 
			12'd2003 :q  <= 20'h4b026; 
			12'd2004 :q  <= 20'h52061; 
			12'd2005 :q  <= 20'h3a061; 
			12'd2006 :q  <= 20'h289ee; 
			12'd2007 :q  <= 20'h1044a; 
			12'd2008 :q  <= 20'h73843; 
			12'd2009 :q  <= 20'h11c63; 
			12'd2010 :q  <= 20'h89063; 
			12'd2011 :q  <= 20'h01063; 
			12'd2012 :q  <= 20'h694c2; 
			12'd2013 :q  <= 20'h24d81; 
			12'd2014 :q  <= 20'h63044; 
			12'd2015 :q  <= 20'h1bc23; 
			12'd2016 :q  <= 20'h5c0c4; 
			12'd2017 :q  <= 20'h1286a; 
			12'd2018 :q  <= 20'h62044; 
			12'd2019 :q  <= 20'h32044; 
			12'd2020 :q  <= 20'h53843; 
			12'd2021 :q  <= 20'h28543; 
			12'd2022 :q  <= 20'h51c62; 
			12'd2023 :q  <= 20'h29922; 
			12'd2024 :q  <= 20'h4a042; 
			12'd2025 :q  <= 20'h12e06; 
			12'd2026 :q  <= 20'h61c42; 
			12'd2027 :q  <= 20'h49443; 
			12'd2028 :q  <= 20'h49c62; 
			12'd2029 :q  <= 20'h2850c; 
			12'd2030 :q  <= 20'h69442; 
			12'd2031 :q  <= 20'h29442; 
			12'd2032 :q  <= 20'h61063; 
			12'd2033 :q  <= 20'h23843; 
			12'd2034 :q  <= 20'h61063; 
			12'd2035 :q  <= 20'h29063; 
			12'd2036 :q  <= 20'h4b846; 
			12'd2037 :q  <= 20'h43862; 
			12'd2038 :q  <= 20'h494c6; 
			12'd2039 :q  <= 20'h294c6; 
			12'd2040 :q  <= 20'h6b422; 
			12'd2041 :q  <= 20'h00942; 
			12'd2042 :q  <= 20'h6b422; 
			12'd2043 :q  <= 20'h29c42; 
			12'd2044 :q  <= 20'h69447; 
			12'd2045 :q  <= 20'h33422; 
			12'd2046 :q  <= 20'h58067; 
			12'd2047 :q  <= 20'h00c50; 
			12'd2048 :q  <= 20'h58067; 
			12'd2049 :q  <= 20'h30067; 
			12'd2050 :q  <= 20'h5c104; 
			12'd2051 :q  <= 20'h0c104; 
			12'd2052 :q  <= 20'h69447; 
			12'd2053 :q  <= 20'h29447; 
			12'd2054 :q  <= 20'h9184e; 
			12'd2055 :q  <= 20'h32864; 
			12'd2056 :q  <= 20'h71c22; 
			12'd2057 :q  <= 20'h00646; 
			12'd2058 :q  <= 20'h71c22; 
			12'd2059 :q  <= 20'h0184e; 
			12'd2060 :q  <= 20'h8806c; 
			12'd2061 :q  <= 20'h01a43; 
			12'd2062 :q  <= 20'h301d0; 
			12'd2063 :q  <= 20'h0006c; 
			12'd2064 :q  <= 20'h68067; 
			12'd2065 :q  <= 20'h29c22; 
			12'd2066 :q  <= 20'h710c6; 
			12'd2067 :q  <= 20'h29ce2; 
			12'd2068 :q  <= 20'h418c9; 
			12'd2069 :q  <= 20'h290c1; 
			12'd2070 :q  <= 20'h680c4; 
			12'd2071 :q  <= 20'h08a4c; 
			12'd2072 :q  <= 20'h18a2c; 
			12'd2073 :q  <= 20'h2b8e3; 
			12'd2074 :q  <= 20'h53823; 
			12'd2075 :q  <= 20'h1b863; 
			12'd2076 :q  <= 20'h710c6; 
			12'd2077 :q  <= 20'h010c6; 
			12'd2078 :q  <= 20'h61483; 
			12'd2079 :q  <= 20'h21483; 
			12'd2080 :q  <= 20'h90046; 
			12'd2081 :q  <= 20'h40489; 
			12'd2082 :q  <= 20'h31902; 
			12'd2083 :q  <= 20'h31482; 
			12'd2084 :q  <= 20'h51443; 
			12'd2085 :q  <= 20'h49423; 
			12'd2086 :q  <= 20'h4a842; 
			12'd2087 :q  <= 20'h02083; 
			12'd2088 :q  <= 20'h30106; 
			12'd2089 :q  <= 20'h080c4; 
			12'd2090 :q  <= 20'h68067; 
			12'd2091 :q  <= 20'h4c042; 
			12'd2092 :q  <= 20'h590ca; 
			12'd2093 :q  <= 20'h02a62; 
			12'd2094 :q  <= 20'h49509; 
			12'd2095 :q  <= 20'h20067; 
			12'd2096 :q  <= 20'h4188c; 
			12'd2097 :q  <= 20'h008c4; 
			12'd2098 :q  <= 20'h43c83; 
			12'd2099 :q  <= 20'h40067; 
			12'd2100 :q  <= 20'h49464; 
			12'd2101 :q  <= 20'h41464; 
			12'd2102 :q  <= 20'h398c1; 
			12'd2103 :q  <= 20'h3b884; 
			12'd2104 :q  <= 20'h6b886; 
			12'd2105 :q  <= 20'h3a028; 
			12'd2106 :q  <= 20'h80048; 
			12'd2107 :q  <= 20'h10048; 
			12'd2108 :q  <= 20'h305c3; 
			12'd2109 :q  <= 20'h3a46a; 
			12'd2110 :q  <= 20'h4b842; 
			12'd2111 :q  <= 20'h39cc8; 
			12'd2112 :q  <= 20'h49c66; 
			12'd2113 :q  <= 20'h3b463; 
			12'd2114 :q  <= 20'h4a442; 
			12'd2115 :q  <= 20'h00642; 
			12'd2116 :q  <= 20'h384ce; 
			12'd2117 :q  <= 20'h0a641; 
			12'd2118 :q  <= 20'h49c42; 
			12'd2119 :q  <= 20'h48c49; 
			12'd2120 :q  <= 20'h93843; 
			12'd2121 :q  <= 20'h3ac61; 
			12'd2122 :q  <= 20'h52064; 
			12'd2123 :q  <= 20'h3b866; 
			12'd2124 :q  <= 20'h52064; 
			12'd2125 :q  <= 20'h3a064; 
			12'd2126 :q  <= 20'h3a4c9; 
			12'd2127 :q  <= 20'h03843; 
			12'd2128 :q  <= 20'h5b022; 
			12'd2129 :q  <= 20'h20d03; 
			12'd2130 :q  <= 20'h01286; 
			12'd2131 :q  <= 20'h4b823; 
			12'd2132 :q  <= 20'h43883; 
			12'd2133 :q  <= 20'h03dc4; 
			12'd2134 :q  <= 20'h0ba46; 
			12'd2135 :q  <= 20'h00146;
			default	 :q  <= 20'h00000;
		endcase	
	end
	assign out = q;
endmodule