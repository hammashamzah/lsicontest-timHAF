module mux_400_to_1_9bit(
	input[8:0] address,
	input[20*20*9 - 1 : 0] image,
	output reg[8:0] out
);
	
		always @(address or image) begin
		case (address)
			9'd0   : out <= image[8 : 0];
			9'd1   : out <= image[17 : 9];
			9'd2   : out <= image[26 : 18];
			9'd3   : out <= image[35 : 27];
			9'd4   : out <= image[44 : 36];
			9'd5   : out <= image[53 : 45];
			9'd6   : out <= image[62 : 54];
			9'd7   : out <= image[71 : 63];
			9'd8   : out <= image[80 : 72];
			9'd9   : out <= image[89 : 81];
			9'd10  : out <= image[98 : 90];
			9'd11  : out <= image[107 : 99];
			9'd12  : out <= image[116 : 108];
			9'd13  : out <= image[125 : 117];
			9'd14  : out <= image[134 : 126];
			9'd15  : out <= image[143 : 135];
			9'd16  : out <= image[152 : 144];
			9'd17  : out <= image[161 : 153];
			9'd18  : out <= image[170 : 162];
			9'd19  : out <= image[179 : 171];
			9'd20  : out <= image[188 : 180];
			9'd21  : out <= image[197 : 189];
			9'd22  : out <= image[206 : 198];
			9'd23  : out <= image[215 : 207];
			9'd24  : out <= image[224 : 216];
			9'd25  : out <= image[233 : 225];
			9'd26  : out <= image[242 : 234];
			9'd27  : out <= image[251 : 243];
			9'd28  : out <= image[260 : 252];
			9'd29  : out <= image[269 : 261];
			9'd30  : out <= image[278 : 270];
			9'd31  : out <= image[287 : 279];
			9'd32  : out <= image[296 : 288];
			9'd33  : out <= image[305 : 297];
			9'd34  : out <= image[314 : 306];
			9'd35  : out <= image[323 : 315];
			9'd36  : out <= image[332 : 324];
			9'd37  : out <= image[341 : 333];
			9'd38  : out <= image[350 : 342];
			9'd39  : out <= image[359 : 351];
			9'd40  : out <= image[368 : 360];
			9'd41  : out <= image[377 : 369];
			9'd42  : out <= image[386 : 378];
			9'd43  : out <= image[395 : 387];
			9'd44  : out <= image[404 : 396];
			9'd45  : out <= image[413 : 405];
			9'd46  : out <= image[422 : 414];
			9'd47  : out <= image[431 : 423];
			9'd48  : out <= image[440 : 432];
			9'd49  : out <= image[449 : 441];
			9'd50  : out <= image[458 : 450];
			9'd51  : out <= image[467 : 459];
			9'd52  : out <= image[476 : 468];
			9'd53  : out <= image[485 : 477];
			9'd54  : out <= image[494 : 486];
			9'd55  : out <= image[503 : 495];
			9'd56  : out <= image[512 : 504];
			9'd57  : out <= image[521 : 513];
			9'd58  : out <= image[530 : 522];
			9'd59  : out <= image[539 : 531];
			9'd60  : out <= image[548 : 540];
			9'd61  : out <= image[557 : 549];
			9'd62  : out <= image[566 : 558];
			9'd63  : out <= image[575 : 567];
			9'd64  : out <= image[584 : 576];
			9'd65  : out <= image[593 : 585];
			9'd66  : out <= image[602 : 594];
			9'd67  : out <= image[611 : 603];
			9'd68  : out <= image[620 : 612];
			9'd69  : out <= image[629 : 621];
			9'd70  : out <= image[638 : 630];
			9'd71  : out <= image[647 : 639];
			9'd72  : out <= image[656 : 648];
			9'd73  : out <= image[665 : 657];
			9'd74  : out <= image[674 : 666];
			9'd75  : out <= image[683 : 675];
			9'd76  : out <= image[692 : 684];
			9'd77  : out <= image[701 : 693];
			9'd78  : out <= image[710 : 702];
			9'd79  : out <= image[719 : 711];
			9'd80  : out <= image[728 : 720];
			9'd81  : out <= image[737 : 729];
			9'd82  : out <= image[746 : 738];
			9'd83  : out <= image[755 : 747];
			9'd84  : out <= image[764 : 756];
			9'd85  : out <= image[773 : 765];
			9'd86  : out <= image[782 : 774];
			9'd87  : out <= image[791 : 783];
			9'd88  : out <= image[800 : 792];
			9'd89  : out <= image[809 : 801];
			9'd90  : out <= image[818 : 810];
			9'd91  : out <= image[827 : 819];
			9'd92  : out <= image[836 : 828];
			9'd93  : out <= image[845 : 837];
			9'd94  : out <= image[854 : 846];
			9'd95  : out <= image[863 : 855];
			9'd96  : out <= image[872 : 864];
			9'd97  : out <= image[881 : 873];
			9'd98  : out <= image[890 : 882];
			9'd99  : out <= image[899 : 891];
			9'd100 : out <= image[908 : 900];
			9'd101 : out <= image[917 : 909];
			9'd102 : out <= image[926 : 918];
			9'd103 : out <= image[935 : 927];
			9'd104 : out <= image[944 : 936];
			9'd105 : out <= image[953 : 945];
			9'd106 : out <= image[962 : 954];
			9'd107 : out <= image[971 : 963];
			9'd108 : out <= image[980 : 972];
			9'd109 : out <= image[989 : 981];
			9'd110 : out <= image[998 : 990];
			9'd111 : out <= image[1007 : 999];
			9'd112 : out <= image[1016 : 1008];
			9'd113 : out <= image[1025 : 1017];
			9'd114 : out <= image[1034 : 1026];
			9'd115 : out <= image[1043 : 1035];
			9'd116 : out <= image[1052 : 1044];
			9'd117 : out <= image[1061 : 1053];
			9'd118 : out <= image[1070 : 1062];
			9'd119 : out <= image[1079 : 1071];
			9'd120 : out <= image[1088 : 1080];
			9'd121 : out <= image[1097 : 1089];
			9'd122 : out <= image[1106 : 1098];
			9'd123 : out <= image[1115 : 1107];
			9'd124 : out <= image[1124 : 1116];
			9'd125 : out <= image[1133 : 1125];
			9'd126 : out <= image[1142 : 1134];
			9'd127 : out <= image[1151 : 1143];
			9'd128 : out <= image[1160 : 1152];
			9'd129 : out <= image[1169 : 1161];
			9'd130 : out <= image[1178 : 1170];
			9'd131 : out <= image[1187 : 1179];
			9'd132 : out <= image[1196 : 1188];
			9'd133 : out <= image[1205 : 1197];
			9'd134 : out <= image[1214 : 1206];
			9'd135 : out <= image[1223 : 1215];
			9'd136 : out <= image[1232 : 1224];
			9'd137 : out <= image[1241 : 1233];
			9'd138 : out <= image[1250 : 1242];
			9'd139 : out <= image[1259 : 1251];
			9'd140 : out <= image[1268 : 1260];
			9'd141 : out <= image[1277 : 1269];
			9'd142 : out <= image[1286 : 1278];
			9'd143 : out <= image[1295 : 1287];
			9'd144 : out <= image[1304 : 1296];
			9'd145 : out <= image[1313 : 1305];
			9'd146 : out <= image[1322 : 1314];
			9'd147 : out <= image[1331 : 1323];
			9'd148 : out <= image[1340 : 1332];
			9'd149 : out <= image[1349 : 1341];
			9'd150 : out <= image[1358 : 1350];
			9'd151 : out <= image[1367 : 1359];
			9'd152 : out <= image[1376 : 1368];
			9'd153 : out <= image[1385 : 1377];
			9'd154 : out <= image[1394 : 1386];
			9'd155 : out <= image[1403 : 1395];
			9'd156 : out <= image[1412 : 1404];
			9'd157 : out <= image[1421 : 1413];
			9'd158 : out <= image[1430 : 1422];
			9'd159 : out <= image[1439 : 1431];
			9'd160 : out <= image[1448 : 1440];
			9'd161 : out <= image[1457 : 1449];
			9'd162 : out <= image[1466 : 1458];
			9'd163 : out <= image[1475 : 1467];
			9'd164 : out <= image[1484 : 1476];
			9'd165 : out <= image[1493 : 1485];
			9'd166 : out <= image[1502 : 1494];
			9'd167 : out <= image[1511 : 1503];
			9'd168 : out <= image[1520 : 1512];
			9'd169 : out <= image[1529 : 1521];
			9'd170 : out <= image[1538 : 1530];
			9'd171 : out <= image[1547 : 1539];
			9'd172 : out <= image[1556 : 1548];
			9'd173 : out <= image[1565 : 1557];
			9'd174 : out <= image[1574 : 1566];
			9'd175 : out <= image[1583 : 1575];
			9'd176 : out <= image[1592 : 1584];
			9'd177 : out <= image[1601 : 1593];
			9'd178 : out <= image[1610 : 1602];
			9'd179 : out <= image[1619 : 1611];
			9'd180 : out <= image[1628 : 1620];
			9'd181 : out <= image[1637 : 1629];
			9'd182 : out <= image[1646 : 1638];
			9'd183 : out <= image[1655 : 1647];
			9'd184 : out <= image[1664 : 1656];
			9'd185 : out <= image[1673 : 1665];
			9'd186 : out <= image[1682 : 1674];
			9'd187 : out <= image[1691 : 1683];
			9'd188 : out <= image[1700 : 1692];
			9'd189 : out <= image[1709 : 1701];
			9'd190 : out <= image[1718 : 1710];
			9'd191 : out <= image[1727 : 1719];
			9'd192 : out <= image[1736 : 1728];
			9'd193 : out <= image[1745 : 1737];
			9'd194 : out <= image[1754 : 1746];
			9'd195 : out <= image[1763 : 1755];
			9'd196 : out <= image[1772 : 1764];
			9'd197 : out <= image[1781 : 1773];
			9'd198 : out <= image[1790 : 1782];
			9'd199 : out <= image[1799 : 1791];
			9'd200 : out <= image[1808 : 1800];
			9'd201 : out <= image[1817 : 1809];
			9'd202 : out <= image[1826 : 1818];
			9'd203 : out <= image[1835 : 1827];
			9'd204 : out <= image[1844 : 1836];
			9'd205 : out <= image[1853 : 1845];
			9'd206 : out <= image[1862 : 1854];
			9'd207 : out <= image[1871 : 1863];
			9'd208 : out <= image[1880 : 1872];
			9'd209 : out <= image[1889 : 1881];
			9'd210 : out <= image[1898 : 1890];
			9'd211 : out <= image[1907 : 1899];
			9'd212 : out <= image[1916 : 1908];
			9'd213 : out <= image[1925 : 1917];
			9'd214 : out <= image[1934 : 1926];
			9'd215 : out <= image[1943 : 1935];
			9'd216 : out <= image[1952 : 1944];
			9'd217 : out <= image[1961 : 1953];
			9'd218 : out <= image[1970 : 1962];
			9'd219 : out <= image[1979 : 1971];
			9'd220 : out <= image[1988 : 1980];
			9'd221 : out <= image[1997 : 1989];
			9'd222 : out <= image[2006 : 1998];
			9'd223 : out <= image[2015 : 2007];
			9'd224 : out <= image[2024 : 2016];
			9'd225 : out <= image[2033 : 2025];
			9'd226 : out <= image[2042 : 2034];
			9'd227 : out <= image[2051 : 2043];
			9'd228 : out <= image[2060 : 2052];
			9'd229 : out <= image[2069 : 2061];
			9'd230 : out <= image[2078 : 2070];
			9'd231 : out <= image[2087 : 2079];
			9'd232 : out <= image[2096 : 2088];
			9'd233 : out <= image[2105 : 2097];
			9'd234 : out <= image[2114 : 2106];
			9'd235 : out <= image[2123 : 2115];
			9'd236 : out <= image[2132 : 2124];
			9'd237 : out <= image[2141 : 2133];
			9'd238 : out <= image[2150 : 2142];
			9'd239 : out <= image[2159 : 2151];
			9'd240 : out <= image[2168 : 2160];
			9'd241 : out <= image[2177 : 2169];
			9'd242 : out <= image[2186 : 2178];
			9'd243 : out <= image[2195 : 2187];
			9'd244 : out <= image[2204 : 2196];
			9'd245 : out <= image[2213 : 2205];
			9'd246 : out <= image[2222 : 2214];
			9'd247 : out <= image[2231 : 2223];
			9'd248 : out <= image[2240 : 2232];
			9'd249 : out <= image[2249 : 2241];
			9'd250 : out <= image[2258 : 2250];
			9'd251 : out <= image[2267 : 2259];
			9'd252 : out <= image[2276 : 2268];
			9'd253 : out <= image[2285 : 2277];
			9'd254 : out <= image[2294 : 2286];
			9'd255 : out <= image[2303 : 2295];
			9'd256 : out <= image[2312 : 2304];
			9'd257 : out <= image[2321 : 2313];
			9'd258 : out <= image[2330 : 2322];
			9'd259 : out <= image[2339 : 2331];
			9'd260 : out <= image[2348 : 2340];
			9'd261 : out <= image[2357 : 2349];
			9'd262 : out <= image[2366 : 2358];
			9'd263 : out <= image[2375 : 2367];
			9'd264 : out <= image[2384 : 2376];
			9'd265 : out <= image[2393 : 2385];
			9'd266 : out <= image[2402 : 2394];
			9'd267 : out <= image[2411 : 2403];
			9'd268 : out <= image[2420 : 2412];
			9'd269 : out <= image[2429 : 2421];
			9'd270 : out <= image[2438 : 2430];
			9'd271 : out <= image[2447 : 2439];
			9'd272 : out <= image[2456 : 2448];
			9'd273 : out <= image[2465 : 2457];
			9'd274 : out <= image[2474 : 2466];
			9'd275 : out <= image[2483 : 2475];
			9'd276 : out <= image[2492 : 2484];
			9'd277 : out <= image[2501 : 2493];
			9'd278 : out <= image[2510 : 2502];
			9'd279 : out <= image[2519 : 2511];
			9'd280 : out <= image[2528 : 2520];
			9'd281 : out <= image[2537 : 2529];
			9'd282 : out <= image[2546 : 2538];
			9'd283 : out <= image[2555 : 2547];
			9'd284 : out <= image[2564 : 2556];
			9'd285 : out <= image[2573 : 2565];
			9'd286 : out <= image[2582 : 2574];
			9'd287 : out <= image[2591 : 2583];
			9'd288 : out <= image[2600 : 2592];
			9'd289 : out <= image[2609 : 2601];
			9'd290 : out <= image[2618 : 2610];
			9'd291 : out <= image[2627 : 2619];
			9'd292 : out <= image[2636 : 2628];
			9'd293 : out <= image[2645 : 2637];
			9'd294 : out <= image[2654 : 2646];
			9'd295 : out <= image[2663 : 2655];
			9'd296 : out <= image[2672 : 2664];
			9'd297 : out <= image[2681 : 2673];
			9'd298 : out <= image[2690 : 2682];
			9'd299 : out <= image[2699 : 2691];
			9'd300 : out <= image[2708 : 2700];
			9'd301 : out <= image[2717 : 2709];
			9'd302 : out <= image[2726 : 2718];
			9'd303 : out <= image[2735 : 2727];
			9'd304 : out <= image[2744 : 2736];
			9'd305 : out <= image[2753 : 2745];
			9'd306 : out <= image[2762 : 2754];
			9'd307 : out <= image[2771 : 2763];
			9'd308 : out <= image[2780 : 2772];
			9'd309 : out <= image[2789 : 2781];
			9'd310 : out <= image[2798 : 2790];
			9'd311 : out <= image[2807 : 2799];
			9'd312 : out <= image[2816 : 2808];
			9'd313 : out <= image[2825 : 2817];
			9'd314 : out <= image[2834 : 2826];
			9'd315 : out <= image[2843 : 2835];
			9'd316 : out <= image[2852 : 2844];
			9'd317 : out <= image[2861 : 2853];
			9'd318 : out <= image[2870 : 2862];
			9'd319 : out <= image[2879 : 2871];
			9'd320 : out <= image[2888 : 2880];
			9'd321 : out <= image[2897 : 2889];
			9'd322 : out <= image[2906 : 2898];
			9'd323 : out <= image[2915 : 2907];
			9'd324 : out <= image[2924 : 2916];
			9'd325 : out <= image[2933 : 2925];
			9'd326 : out <= image[2942 : 2934];
			9'd327 : out <= image[2951 : 2943];
			9'd328 : out <= image[2960 : 2952];
			9'd329 : out <= image[2969 : 2961];
			9'd330 : out <= image[2978 : 2970];
			9'd331 : out <= image[2987 : 2979];
			9'd332 : out <= image[2996 : 2988];
			9'd333 : out <= image[3005 : 2997];
			9'd334 : out <= image[3014 : 3006];
			9'd335 : out <= image[3023 : 3015];
			9'd336 : out <= image[3032 : 3024];
			9'd337 : out <= image[3041 : 3033];
			9'd338 : out <= image[3050 : 3042];
			9'd339 : out <= image[3059 : 3051];
			9'd340 : out <= image[3068 : 3060];
			9'd341 : out <= image[3077 : 3069];
			9'd342 : out <= image[3086 : 3078];
			9'd343 : out <= image[3095 : 3087];
			9'd344 : out <= image[3104 : 3096];
			9'd345 : out <= image[3113 : 3105];
			9'd346 : out <= image[3122 : 3114];
			9'd347 : out <= image[3131 : 3123];
			9'd348 : out <= image[3140 : 3132];
			9'd349 : out <= image[3149 : 3141];
			9'd350 : out <= image[3158 : 3150];
			9'd351 : out <= image[3167 : 3159];
			9'd352 : out <= image[3176 : 3168];
			9'd353 : out <= image[3185 : 3177];
			9'd354 : out <= image[3194 : 3186];
			9'd355 : out <= image[3203 : 3195];
			9'd356 : out <= image[3212 : 3204];
			9'd357 : out <= image[3221 : 3213];
			9'd358 : out <= image[3230 : 3222];
			9'd359 : out <= image[3239 : 3231];
			9'd360 : out <= image[3248 : 3240];
			9'd361 : out <= image[3257 : 3249];
			9'd362 : out <= image[3266 : 3258];
			9'd363 : out <= image[3275 : 3267];
			9'd364 : out <= image[3284 : 3276];
			9'd365 : out <= image[3293 : 3285];
			9'd366 : out <= image[3302 : 3294];
			9'd367 : out <= image[3311 : 3303];
			9'd368 : out <= image[3320 : 3312];
			9'd369 : out <= image[3329 : 3321];
			9'd370 : out <= image[3338 : 3330];
			9'd371 : out <= image[3347 : 3339];
			9'd372 : out <= image[3356 : 3348];
			9'd373 : out <= image[3365 : 3357];
			9'd374 : out <= image[3374 : 3366];
			9'd375 : out <= image[3383 : 3375];
			9'd376 : out <= image[3392 : 3384];
			9'd377 : out <= image[3401 : 3393];
			9'd378 : out <= image[3410 : 3402];
			9'd379 : out <= image[3419 : 3411];
			9'd380 : out <= image[3428 : 3420];
			9'd381 : out <= image[3437 : 3429];
			9'd382 : out <= image[3446 : 3438];
			9'd383 : out <= image[3455 : 3447];
			9'd384 : out <= image[3464 : 3456];
			9'd385 : out <= image[3473 : 3465];
			9'd386 : out <= image[3482 : 3474];
			9'd387 : out <= image[3491 : 3483];
			9'd388 : out <= image[3500 : 3492];
			9'd389 : out <= image[3509 : 3501];
			9'd390 : out <= image[3518 : 3510];
			9'd391 : out <= image[3527 : 3519];
			9'd392 : out <= image[3536 : 3528];
			9'd393 : out <= image[3545 : 3537];
			9'd394 : out <= image[3554 : 3546];
			9'd395 : out <= image[3563 : 3555];
			9'd396 : out <= image[3572 : 3564];
			9'd397 : out <= image[3581 : 3573];
			9'd398 : out <= image[3590 : 3582];
			9'd399 : out <= image[3599 : 3591];
			default : out <= 9'b000000000;
		endcase
	end
endmodule