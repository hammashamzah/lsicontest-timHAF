`define n WindowSize

module IntegralBuffer
(

);


endmodule 