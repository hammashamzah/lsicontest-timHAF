module rect3_rom(
	input [11:0] addr,
	input clk,
	output[22:0] out
);
	reg[22:0] q;

	always @(posedge clk)
	begin
		case(addr)
			12'd1    : q <= 23'h000000;
			12'd2    : q <= 23'h000000;
			12'd3    : q <= 23'h000000;
			12'd4    : q <= 23'h000000;
			12'd5    : q <= 23'h000000;
			12'd6    : q <= 23'h000000;
			12'd7    : q <= 23'h000000;
			12'd8    : q <= 23'h000000;
			12'd9    : q <= 23'h000000;
			12'd10   : q <= 23'h000000;
			12'd11   : q <= 23'h000000;
			12'd12   : q <= 23'h000000;
			12'd13   : q <= 23'h000000;
			12'd14   : q <= 23'h000000;
			12'd15   : q <= 23'h000000;
			12'd16   : q <= 23'h231846;
			12'd17   : q <= 23'h000000;
			12'd18   : q <= 23'h000000;
			12'd19   : q <= 23'h000000;
			12'd20   : q <= 23'h000000;
			12'd21   : q <= 23'h000000;
			12'd22   : q <= 23'h000000;
			12'd23   : q <= 23'h000000;
			12'd24   : q <= 23'h000000;
			12'd25   : q <= 23'h000000;
			12'd26   : q <= 23'h000000;
			12'd27   : q <= 23'h000000;
			12'd28   : q <= 23'h000000;
			12'd29   : q <= 23'h000000;
			12'd30   : q <= 23'h000000;
			12'd31   : q <= 23'h000000;
			12'd32   : q <= 23'h24a524;
			12'd33   : q <= 23'h2444a2;
			12'd34   : q <= 23'h229444;
			12'd35   : q <= 23'h21ace5;
			12'd36   : q <= 23'h000000;
			12'd37   : q <= 23'h000000;
			12'd38   : q <= 23'h000000;
			12'd39   : q <= 23'h000000;
			12'd40   : q <= 23'h000000;
			12'd41   : q <= 23'h000000;
			12'd42   : q <= 23'h000000;
			12'd43   : q <= 23'h000000;
			12'd44   : q <= 23'h000000;
			12'd45   : q <= 23'h000000;
			12'd46   : q <= 23'h259883;
			12'd47   : q <= 23'h000000;
			12'd48   : q <= 23'h000000;
			12'd49   : q <= 23'h000000;
			12'd50   : q <= 23'h2444a2;
			12'd51   : q <= 23'h000000;
			12'd52   : q <= 23'h000000;
			12'd53   : q <= 23'h000000;
			12'd54   : q <= 23'h2224c5;
			12'd55   : q <= 23'h000000;
			12'd56   : q <= 23'h000000;
			12'd57   : q <= 23'h000000;
			12'd58   : q <= 23'h000000;
			12'd59   : q <= 23'h234462;
			12'd60   : q <= 23'h000000;
			12'd61   : q <= 23'h000000;
			12'd62   : q <= 23'h000000;
			12'd63   : q <= 23'h000000;
			12'd64   : q <= 23'h000000;
			12'd65   : q <= 23'h000000;
			12'd66   : q <= 23'h000000;
			12'd67   : q <= 23'h000000;
			12'd68   : q <= 23'h000000;
			12'd69   : q <= 23'h000000;
			12'd70   : q <= 23'h000000;
			12'd71   : q <= 23'h000000;
			12'd72   : q <= 23'h000000;
			12'd73   : q <= 23'h000000;
			12'd74   : q <= 23'h000000;
			12'd75   : q <= 23'h000000;
			12'd76   : q <= 23'h20b122;
			12'd77   : q <= 23'h000000;
			12'd78   : q <= 23'h000000;
			12'd79   : q <= 23'h000000;
			12'd80   : q <= 23'h000000;
			12'd81   : q <= 23'h000000;
			12'd82   : q <= 23'h000000;
			12'd83   : q <= 23'h000000;
			12'd84   : q <= 23'h000000;
			12'd85   : q <= 23'h000000;
			12'd86   : q <= 23'h000000;
			12'd87   : q <= 23'h000000;
			12'd88   : q <= 23'h000000;
			12'd89   : q <= 23'h000000;
			12'd90   : q <= 23'h000000;
			12'd91   : q <= 23'h000000;
			12'd92   : q <= 23'h000000;
			12'd93   : q <= 23'h248842;
			12'd94   : q <= 23'h000000;
			12'd95   : q <= 23'h000000;
			12'd96   : q <= 23'h000000;
			12'd97   : q <= 23'h000000;
			12'd98   : q <= 23'h000000;
			12'd99   : q <= 23'h000000;
			12'd100  : q <= 23'h000000; 
			12'd101  : q <= 23'h000000; 
			12'd102  : q <= 23'h000000; 
			12'd103  : q <= 23'h000000; 
			12'd104  : q <= 23'h000000; 
			12'd105  : q <= 23'h000000; 
			12'd106  : q <= 23'h000000; 
			12'd107  : q <= 23'h240842; 
			12'd108  : q <= 23'h000000; 
			12'd109  : q <= 23'h000000; 
			12'd110  : q <= 23'h2528a6; 
			12'd111  : q <= 23'h000000; 
			12'd112  : q <= 23'h2424c7; 
			12'd113  : q <= 23'h000000; 
			12'd114  : q <= 23'h000000; 
			12'd115  : q <= 23'h000000; 
			12'd116  : q <= 23'h000000; 
			12'd117  : q <= 23'h000000; 
			12'd118  : q <= 23'h000000; 
			12'd119  : q <= 23'h231c65; 
			12'd120  : q <= 23'h000000; 
			12'd121  : q <= 23'h23c483; 
			12'd122  : q <= 23'h000000; 
			12'd123  : q <= 23'h000000; 
			12'd124  : q <= 23'h000000; 
			12'd125  : q <= 23'h24b0e3; 
			12'd126  : q <= 23'h000000; 
			12'd127  : q <= 23'h253484; 
			12'd128  : q <= 23'h000000; 
			12'd129  : q <= 23'h000000; 
			12'd130  : q <= 23'h000000; 
			12'd131  : q <= 23'h000000; 
			12'd132  : q <= 23'h212524; 
			12'd133  : q <= 23'h000000; 
			12'd134  : q <= 23'h000000; 
			12'd135  : q <= 23'h000000; 
			12'd136  : q <= 23'h000000; 
			12'd137  : q <= 23'h000000; 
			12'd138  : q <= 23'h242886; 
			12'd139  : q <= 23'h000000; 
			12'd140  : q <= 23'h000000; 
			12'd141  : q <= 23'h000000; 
			12'd142  : q <= 23'h000000; 
			12'd143  : q <= 23'h000000; 
			12'd144  : q <= 23'h000000; 
			12'd145  : q <= 23'h000000; 
			12'd146  : q <= 23'h000000; 
			12'd147  : q <= 23'h000000; 
			12'd148  : q <= 23'h2234c6; 
			12'd149  : q <= 23'h000000; 
			12'd150  : q <= 23'h000000; 
			12'd151  : q <= 23'h000000; 
			12'd152  : q <= 23'h000000; 
			12'd153  : q <= 23'h000000; 
			12'd154  : q <= 23'h000000; 
			12'd155  : q <= 23'h000000; 
			12'd156  : q <= 23'h000000; 
			12'd157  : q <= 23'h000000; 
			12'd158  : q <= 23'h000000; 
			12'd159  : q <= 23'h000000; 
			12'd160  : q <= 23'h000000; 
			12'd161  : q <= 23'h000000; 
			12'd162  : q <= 23'h000000; 
			12'd163  : q <= 23'h000000; 
			12'd164  : q <= 23'h000000; 
			12'd165  : q <= 23'h000000; 
			12'd166  : q <= 23'h000000; 
			12'd167  : q <= 23'h000000; 
			12'd168  : q <= 23'h000000; 
			12'd169  : q <= 23'h24b085; 
			12'd170  : q <= 23'h2228c6; 
			12'd171  : q <= 23'h000000; 
			12'd172  : q <= 23'h000000; 
			12'd173  : q <= 23'h000000; 
			12'd174  : q <= 23'h000000; 
			12'd175  : q <= 23'h000000; 
			12'd176  : q <= 23'h000000; 
			12'd177  : q <= 23'h000000; 
			12'd178  : q <= 23'h000000; 
			12'd179  : q <= 23'h000000; 
			12'd180  : q <= 23'h000000; 
			12'd181  : q <= 23'h000000; 
			12'd182  : q <= 23'h000000; 
			12'd183  : q <= 23'h229844; 
			12'd184  : q <= 23'h000000; 
			12'd185  : q <= 23'h000000; 
			12'd186  : q <= 23'h000000; 
			12'd187  : q <= 23'h000000; 
			12'd188  : q <= 23'h000000; 
			12'd189  : q <= 23'h000000; 
			12'd190  : q <= 23'h000000; 
			12'd191  : q <= 23'h000000; 
			12'd192  : q <= 23'h203143; 
			12'd193  : q <= 23'h000000; 
			12'd194  : q <= 23'h000000; 
			12'd195  : q <= 23'h000000; 
			12'd196  : q <= 23'h000000; 
			12'd197  : q <= 23'h000000; 
			12'd198  : q <= 23'h000000; 
			12'd199  : q <= 23'h000000; 
			12'd200  : q <= 23'h2324e2; 
			12'd201  : q <= 23'h000000; 
			12'd202  : q <= 23'h000000; 
			12'd203  : q <= 23'h000000; 
			12'd204  : q <= 23'h22b4c4; 
			12'd205  : q <= 23'h000000; 
			12'd206  : q <= 23'h000000; 
			12'd207  : q <= 23'h000000; 
			12'd208  : q <= 23'h261863; 
			12'd209  : q <= 23'h000000; 
			12'd210  : q <= 23'h242887; 
			12'd211  : q <= 23'h000000; 
			12'd212  : q <= 23'h261864; 
			12'd213  : q <= 23'h229864; 
			12'd214  : q <= 23'h000000; 
			12'd215  : q <= 23'h242887; 
			12'd216  : q <= 23'h000000; 
			12'd217  : q <= 23'h000000; 
			12'd218  : q <= 23'h000000; 
			12'd219  : q <= 23'h000000; 
			12'd220  : q <= 23'h000000; 
			12'd221  : q <= 23'h000000; 
			12'd222  : q <= 23'h000000; 
			12'd223  : q <= 23'h000000; 
			12'd224  : q <= 23'h000000; 
			12'd225  : q <= 23'h253502; 
			12'd226  : q <= 23'h26a462; 
			12'd227  : q <= 23'h000000; 
			12'd228  : q <= 23'h000000; 
			12'd229  : q <= 23'h000000; 
			12'd230  : q <= 23'h000000; 
			12'd231  : q <= 23'h000000; 
			12'd232  : q <= 23'h000000; 
			12'd233  : q <= 23'h000000; 
			12'd234  : q <= 23'h000000; 
			12'd235  : q <= 23'h000000; 
			12'd236  : q <= 23'h000000; 
			12'd237  : q <= 23'h000000; 
			12'd238  : q <= 23'h000000; 
			12'd239  : q <= 23'h000000; 
			12'd240  : q <= 23'h2228c3; 
			12'd241  : q <= 23'h000000; 
			12'd242  : q <= 23'h000000; 
			12'd243  : q <= 23'h000000; 
			12'd244  : q <= 23'h000000; 
			12'd245  : q <= 23'h000000; 
			12'd246  : q <= 23'h000000; 
			12'd247  : q <= 23'h000000; 
			12'd248  : q <= 23'h000000; 
			12'd249  : q <= 23'h22a4a2; 
			12'd250  : q <= 23'h000000; 
			12'd251  : q <= 23'h000000; 
			12'd252  : q <= 23'h000000; 
			12'd253  : q <= 23'h000000; 
			12'd254  : q <= 23'h254842; 
			12'd255  : q <= 23'h000000; 
			12'd256  : q <= 23'h000000; 
			12'd257  : q <= 23'h000000; 
			12'd258  : q <= 23'h000000; 
			12'd259  : q <= 23'h000000; 
			12'd260  : q <= 23'h000000; 
			12'd261  : q <= 23'h000000; 
			12'd262  : q <= 23'h000000; 
			12'd263  : q <= 23'h000000; 
			12'd264  : q <= 23'h000000; 
			12'd265  : q <= 23'h000000; 
			12'd266  : q <= 23'h000000; 
			12'd267  : q <= 23'h000000; 
			12'd268  : q <= 23'h000000; 
			12'd269  : q <= 23'h000000; 
			12'd270  : q <= 23'h000000; 
			12'd271  : q <= 23'h000000; 
			12'd272  : q <= 23'h000000; 
			12'd273  : q <= 23'h000000; 
			12'd274  : q <= 23'h000000; 
			12'd275  : q <= 23'h000000; 
			12'd276  : q <= 23'h000000; 
			12'd277  : q <= 23'h000000; 
			12'd278  : q <= 23'h000000; 
			12'd279  : q <= 23'h000000; 
			12'd280  : q <= 23'h000000; 
			12'd281  : q <= 23'h26a461; 
			12'd282  : q <= 23'h000000; 
			12'd283  : q <= 23'h203d42; 
			12'd284  : q <= 23'h000000; 
			12'd285  : q <= 23'h000000; 
			12'd286  : q <= 23'h222461; 
			12'd287  : q <= 23'h200d41; 
			12'd288  : q <= 23'h000000; 
			12'd289  : q <= 23'h23c063; 
			12'd290  : q <= 23'h000000; 
			12'd291  : q <= 23'h000000; 
			12'd292  : q <= 23'h000000; 
			12'd293  : q <= 23'h2228e6; 
			12'd294  : q <= 23'h000000; 
			12'd295  : q <= 23'h000000; 
			12'd296  : q <= 23'h000000; 
			12'd297  : q <= 23'h000000; 
			12'd298  : q <= 23'h229845; 
			12'd299  : q <= 23'h000000; 
			12'd300  : q <= 23'h000000; 
			12'd301  : q <= 23'h000000; 
			12'd302  : q <= 23'h000000; 
			12'd303  : q <= 23'h000000; 
			12'd304  : q <= 23'h252cc6; 
			12'd305  : q <= 23'h000000; 
			12'd306  : q <= 23'h000000; 
			12'd307  : q <= 23'h218ce1; 
			12'd308  : q <= 23'h000000; 
			12'd309  : q <= 23'h000000; 
			12'd310  : q <= 23'h000000; 
			12'd311  : q <= 23'h000000; 
			12'd312  : q <= 23'h000000; 
			12'd313  : q <= 23'h000000; 
			12'd314  : q <= 23'h000000; 
			12'd315  : q <= 23'h000000; 
			12'd316  : q <= 23'h000000; 
			12'd317  : q <= 23'h000000; 
			12'd318  : q <= 23'h000000; 
			12'd319  : q <= 23'h000000; 
			12'd320  : q <= 23'h000000; 
			12'd321  : q <= 23'h000000; 
			12'd322  : q <= 23'h000000; 
			12'd323  : q <= 23'h201543; 
			12'd324  : q <= 23'h231c65; 
			12'd325  : q <= 23'h000000; 
			12'd326  : q <= 23'h000000; 
			12'd327  : q <= 23'h000000; 
			12'd328  : q <= 23'h000000; 
			12'd329  : q <= 23'h000000; 
			12'd330  : q <= 23'h234043; 
			12'd331  : q <= 23'h231886; 
			12'd332  : q <= 23'h000000; 
			12'd333  : q <= 23'h000000; 
			12'd334  : q <= 23'h000000; 
			12'd335  : q <= 23'h000000; 
			12'd336  : q <= 23'h000000; 
			12'd337  : q <= 23'h000000; 
			12'd338  : q <= 23'h000000; 
			12'd339  : q <= 23'h000000; 
			12'd340  : q <= 23'h000000; 
			12'd341  : q <= 23'h000000; 
			12'd342  : q <= 23'h000000; 
			12'd343  : q <= 23'h000000; 
			12'd344  : q <= 23'h000000; 
			12'd345  : q <= 23'h000000; 
			12'd346  : q <= 23'h000000; 
			12'd347  : q <= 23'h000000; 
			12'd348  : q <= 23'h000000; 
			12'd349  : q <= 23'h000000; 
			12'd350  : q <= 23'h000000; 
			12'd351  : q <= 23'h000000; 
			12'd352  : q <= 23'h000000; 
			12'd353  : q <= 23'h000000; 
			12'd354  : q <= 23'h000000; 
			12'd355  : q <= 23'h000000; 
			12'd356  : q <= 23'h000000; 
			12'd357  : q <= 23'h000000; 
			12'd358  : q <= 23'h000000; 
			12'd359  : q <= 23'h000000; 
			12'd360  : q <= 23'h000000; 
			12'd361  : q <= 23'h000000; 
			12'd362  : q <= 23'h000000; 
			12'd363  : q <= 23'h000000; 
			12'd364  : q <= 23'h000000; 
			12'd365  : q <= 23'h000000; 
			12'd366  : q <= 23'h2544e2; 
			12'd367  : q <= 23'h211102; 
			12'd368  : q <= 23'h000000; 
			12'd369  : q <= 23'h000000; 
			12'd370  : q <= 23'h000000; 
			12'd371  : q <= 23'h26a462; 
			12'd372  : q <= 23'h000000; 
			12'd373  : q <= 23'h26a462; 
			12'd374  : q <= 23'h222462; 
			12'd375  : q <= 23'h000000; 
			12'd376  : q <= 23'h000000; 
			12'd377  : q <= 23'h000000; 
			12'd378  : q <= 23'h000000; 
			12'd379  : q <= 23'h000000; 
			12'd380  : q <= 23'h231022; 
			12'd381  : q <= 23'h000000; 
			12'd382  : q <= 23'h000000; 
			12'd383  : q <= 23'h000000; 
			12'd384  : q <= 23'h000000; 
			12'd385  : q <= 23'h000000; 
			12'd386  : q <= 23'h24a865; 
			12'd387  : q <= 23'h24ac86; 
			12'd388  : q <= 23'h000000; 
			12'd389  : q <= 23'h000000; 
			12'd390  : q <= 23'h000000; 
			12'd391  : q <= 23'h000000; 
			12'd392  : q <= 23'h000000; 
			12'd393  : q <= 23'h000000; 
			12'd394  : q <= 23'h000000; 
			12'd395  : q <= 23'h000000; 
			12'd396  : q <= 23'h000000; 
			12'd397  : q <= 23'h000000; 
			12'd398  : q <= 23'h000000; 
			12'd399  : q <= 23'h000000; 
			12'd400  : q <= 23'h000000; 
			12'd401  : q <= 23'h000000; 
			12'd402  : q <= 23'h23c063; 
			12'd403  : q <= 23'h000000; 
			12'd404  : q <= 23'h000000; 
			12'd405  : q <= 23'h000000; 
			12'd406  : q <= 23'h000000; 
			12'd407  : q <= 23'h000000; 
			12'd408  : q <= 23'h000000; 
			12'd409  : q <= 23'h000000; 
			12'd410  : q <= 23'h000000; 
			12'd411  : q <= 23'h000000; 
			12'd412  : q <= 23'h000000; 
			12'd413  : q <= 23'h000000; 
			12'd414  : q <= 23'h000000; 
			12'd415  : q <= 23'h000000; 
			12'd416  : q <= 23'h000000; 
			12'd417  : q <= 23'h000000; 
			12'd418  : q <= 23'h000000; 
			12'd419  : q <= 23'h000000; 
			12'd420  : q <= 23'h210d22; 
			12'd421  : q <= 23'h000000; 
			12'd422  : q <= 23'h2294a3; 
			12'd423  : q <= 23'h000000; 
			12'd424  : q <= 23'h000000; 
			12'd425  : q <= 23'h000000; 
			12'd426  : q <= 23'h000000; 
			12'd427  : q <= 23'h000000; 
			12'd428  : q <= 23'h000000; 
			12'd429  : q <= 23'h000000; 
			12'd430  : q <= 23'h000000; 
			12'd431  : q <= 23'h000000; 
			12'd432  : q <= 23'h000000; 
			12'd433  : q <= 23'h000000; 
			12'd434  : q <= 23'h000000; 
			12'd435  : q <= 23'h000000; 
			12'd436  : q <= 23'h000000; 
			12'd437  : q <= 23'h000000; 
			12'd438  : q <= 23'h000000; 
			12'd439  : q <= 23'h000000; 
			12'd440  : q <= 23'h000000; 
			12'd441  : q <= 23'h000000; 
			12'd442  : q <= 23'h000000; 
			12'd443  : q <= 23'h22c443; 
			12'd444  : q <= 23'h000000; 
			12'd445  : q <= 23'h000000; 
			12'd446  : q <= 23'h000000; 
			12'd447  : q <= 23'h000000; 
			12'd448  : q <= 23'h000000; 
			12'd449  : q <= 23'h000000; 
			12'd450  : q <= 23'h000000; 
			12'd451  : q <= 23'h000000; 
			12'd452  : q <= 23'h000000; 
			12'd453  : q <= 23'h000000; 
			12'd454  : q <= 23'h000000; 
			12'd455  : q <= 23'h000000; 
			12'd456  : q <= 23'h000000; 
			12'd457  : q <= 23'h239c21; 
			12'd458  : q <= 23'h213522; 
			12'd459  : q <= 23'h239c21; 
			12'd460  : q <= 23'h000000; 
			12'd461  : q <= 23'h000000; 
			12'd462  : q <= 23'h000000; 
			12'd463  : q <= 23'h000000; 
			12'd464  : q <= 23'h000000; 
			12'd465  : q <= 23'h000000; 
			12'd466  : q <= 23'h24a462; 
			12'd467  : q <= 23'h000000; 
			12'd468  : q <= 23'h25c442; 
			12'd469  : q <= 23'h000000; 
			12'd470  : q <= 23'h000000; 
			12'd471  : q <= 23'h23c442; 
			12'd472  : q <= 23'h000000; 
			12'd473  : q <= 23'h000000; 
			12'd474  : q <= 23'h000000; 
			12'd475  : q <= 23'h000000; 
			12'd476  : q <= 23'h000000; 
			12'd477  : q <= 23'h000000; 
			12'd478  : q <= 23'h000000; 
			12'd479  : q <= 23'h000000; 
			12'd480  : q <= 23'h000000; 
			12'd481  : q <= 23'h000000; 
			12'd482  : q <= 23'h000000; 
			12'd483  : q <= 23'h000000; 
			12'd484  : q <= 23'h000000; 
			12'd485  : q <= 23'h000000; 
			12'd486  : q <= 23'h000000; 
			12'd487  : q <= 23'h000000; 
			12'd488  : q <= 23'h000000; 
			12'd489  : q <= 23'h000000; 
			12'd490  : q <= 23'h000000; 
			12'd491  : q <= 23'h000000; 
			12'd492  : q <= 23'h000000; 
			12'd493  : q <= 23'h000000; 
			12'd494  : q <= 23'h000000; 
			12'd495  : q <= 23'h000000; 
			12'd496  : q <= 23'h21c0e2; 
			12'd497  : q <= 23'h24c061; 
			12'd498  : q <= 23'h000000; 
			12'd499  : q <= 23'h000000; 
			12'd500  : q <= 23'h000000; 
			12'd501  : q <= 23'h000000; 
			12'd502  : q <= 23'h000000; 
			12'd503  : q <= 23'h000000; 
			12'd504  : q <= 23'h000000; 
			12'd505  : q <= 23'h000000; 
			12'd506  : q <= 23'h000000; 
			12'd507  : q <= 23'h000000; 
			12'd508  : q <= 23'h000000; 
			12'd509  : q <= 23'h000000; 
			12'd510  : q <= 23'h000000; 
			12'd511  : q <= 23'h2528e4; 
			12'd512  : q <= 23'h000000; 
			12'd513  : q <= 23'h24a8c6; 
			12'd514  : q <= 23'h000000; 
			12'd515  : q <= 23'h000000; 
			12'd516  : q <= 23'h000000; 
			12'd517  : q <= 23'h000000; 
			12'd518  : q <= 23'h000000; 
			12'd519  : q <= 23'h000000; 
			12'd520  : q <= 23'h000000; 
			12'd521  : q <= 23'h241c61; 
			12'd522  : q <= 23'h000000; 
			12'd523  : q <= 23'h000000; 
			12'd524  : q <= 23'h000000; 
			12'd525  : q <= 23'h24b502; 
			12'd526  : q <= 23'h000000; 
			12'd527  : q <= 23'h000000; 
			12'd528  : q <= 23'h000000; 
			12'd529  : q <= 23'h000000; 
			12'd530  : q <= 23'h000000; 
			12'd531  : q <= 23'h000000; 
			12'd532  : q <= 23'h000000; 
			12'd533  : q <= 23'h000000; 
			12'd534  : q <= 23'h000000; 
			12'd535  : q <= 23'h000000; 
			12'd536  : q <= 23'h000000; 
			12'd537  : q <= 23'h000000; 
			12'd538  : q <= 23'h000000; 
			12'd539  : q <= 23'h000000; 
			12'd540  : q <= 23'h000000; 
			12'd541  : q <= 23'h000000; 
			12'd542  : q <= 23'h000000; 
			12'd543  : q <= 23'h000000; 
			12'd544  : q <= 23'h000000; 
			12'd545  : q <= 23'h000000; 
			12'd546  : q <= 23'h000000; 
			12'd547  : q <= 23'h000000; 
			12'd548  : q <= 23'h000000; 
			12'd549  : q <= 23'h000000; 
			12'd550  : q <= 23'h000000; 
			12'd551  : q <= 23'h252907; 
			12'd552  : q <= 23'h282c49; 
			12'd553  : q <= 23'h000000; 
			12'd554  : q <= 23'h282c49; 
			12'd555  : q <= 23'h000000; 
			12'd556  : q <= 23'h000000; 
			12'd557  : q <= 23'h000000; 
			12'd558  : q <= 23'h000000; 
			12'd559  : q <= 23'h000000; 
			12'd560  : q <= 23'h000000; 
			12'd561  : q <= 23'h000000; 
			12'd562  : q <= 23'h000000; 
			12'd563  : q <= 23'h000000; 
			12'd564  : q <= 23'h000000; 
			12'd565  : q <= 23'h000000; 
			12'd566  : q <= 23'h22a4a4; 
			12'd567  : q <= 23'h2524c2; 
			12'd568  : q <= 23'h000000; 
			12'd569  : q <= 23'h24a462; 
			12'd570  : q <= 23'h000000; 
			12'd571  : q <= 23'h24c862; 
			12'd572  : q <= 23'h000000; 
			12'd573  : q <= 23'h000000; 
			12'd574  : q <= 23'h000000; 
			12'd575  : q <= 23'h000000; 
			12'd576  : q <= 23'h000000; 
			12'd577  : q <= 23'h000000; 
			12'd578  : q <= 23'h000000; 
			12'd579  : q <= 23'h000000; 
			12'd580  : q <= 23'h000000; 
			12'd581  : q <= 23'h000000; 
			12'd582  : q <= 23'h000000; 
			12'd583  : q <= 23'h000000; 
			12'd584  : q <= 23'h000000; 
			12'd585  : q <= 23'h000000; 
			12'd586  : q <= 23'h000000; 
			12'd587  : q <= 23'h000000; 
			12'd588  : q <= 23'h000000; 
			12'd589  : q <= 23'h000000; 
			12'd590  : q <= 23'h000000; 
			12'd591  : q <= 23'h000000; 
			12'd592  : q <= 23'h000000; 
			12'd593  : q <= 23'h000000; 
			12'd594  : q <= 23'h000000; 
			12'd595  : q <= 23'h000000; 
			12'd596  : q <= 23'h000000; 
			12'd597  : q <= 23'h000000; 
			12'd598  : q <= 23'h000000; 
			12'd599  : q <= 23'h000000; 
			12'd600  : q <= 23'h000000; 
			12'd601  : q <= 23'h25ac21; 
			12'd602  : q <= 23'h000000; 
			12'd603  : q <= 23'h000000; 
			12'd604  : q <= 23'h000000; 
			12'd605  : q <= 23'h000000; 
			12'd606  : q <= 23'h000000; 
			12'd607  : q <= 23'h25ac21; 
			12'd608  : q <= 23'h000000; 
			12'd609  : q <= 23'h000000; 
			12'd610  : q <= 23'h000000; 
			12'd611  : q <= 23'h000000; 
			12'd612  : q <= 23'h000000; 
			12'd613  : q <= 23'h000000; 
			12'd614  : q <= 23'h000000; 
			12'd615  : q <= 23'h000000; 
			12'd616  : q <= 23'h219865; 
			12'd617  : q <= 23'h000000; 
			12'd618  : q <= 23'h000000; 
			12'd619  : q <= 23'h000000; 
			12'd620  : q <= 23'h000000; 
			12'd621  : q <= 23'h000000; 
			12'd622  : q <= 23'h000000; 
			12'd623  : q <= 23'h25ac21; 
			12'd624  : q <= 23'h242c21; 
			12'd625  : q <= 23'h000000; 
			12'd626  : q <= 23'h000000; 
			12'd627  : q <= 23'h000000; 
			12'd628  : q <= 23'h000000; 
			12'd629  : q <= 23'h22b0a5; 
			12'd630  : q <= 23'h23cc81; 
			12'd631  : q <= 23'h000000; 
			12'd632  : q <= 23'h000000; 
			12'd633  : q <= 23'h000000; 
			12'd634  : q <= 23'h000000; 
			12'd635  : q <= 23'h000000; 
			12'd636  : q <= 23'h244021; 
			12'd637  : q <= 23'h000000; 
			12'd638  : q <= 23'h000000; 
			12'd639  : q <= 23'h000000; 
			12'd640  : q <= 23'h000000; 
			12'd641  : q <= 23'h000000; 
			12'd642  : q <= 23'h000000; 
			12'd643  : q <= 23'h000000; 
			12'd644  : q <= 23'h000000; 
			12'd645  : q <= 23'h000000; 
			12'd646  : q <= 23'h000000; 
			12'd647  : q <= 23'h000000; 
			12'd648  : q <= 23'h000000; 
			12'd649  : q <= 23'h000000; 
			12'd650  : q <= 23'h000000; 
			12'd651  : q <= 23'h000000; 
			12'd652  : q <= 23'h24b025; 
			12'd653  : q <= 23'h000000; 
			12'd654  : q <= 23'h000000; 
			12'd655  : q <= 23'h000000; 
			12'd656  : q <= 23'h000000; 
			12'd657  : q <= 23'h000000; 
			12'd658  : q <= 23'h000000; 
			12'd659  : q <= 23'h000000; 
			12'd660  : q <= 23'h000000; 
			12'd661  : q <= 23'h000000; 
			12'd662  : q <= 23'h000000; 
			12'd663  : q <= 23'h000000; 
			12'd664  : q <= 23'h000000; 
			12'd665  : q <= 23'h000000; 
			12'd666  : q <= 23'h000000; 
			12'd667  : q <= 23'h292829; 
			12'd668  : q <= 23'h000000; 
			12'd669  : q <= 23'h292829; 
			12'd670  : q <= 23'h21c443; 
			12'd671  : q <= 23'h000000; 
			12'd672  : q <= 23'h21bc65; 
			12'd673  : q <= 23'h000000; 
			12'd674  : q <= 23'h000000; 
			12'd675  : q <= 23'h000000; 
			12'd676  : q <= 23'h252923; 
			12'd677  : q <= 23'h000000; 
			12'd678  : q <= 23'h000000; 
			12'd679  : q <= 23'h000000; 
			12'd680  : q <= 23'h000000; 
			12'd681  : q <= 23'h000000; 
			12'd682  : q <= 23'h000000; 
			12'd683  : q <= 23'h000000; 
			12'd684  : q <= 23'h26a442; 
			12'd685  : q <= 23'h22a442; 
			12'd686  : q <= 23'h000000; 
			12'd687  : q <= 23'h000000; 
			12'd688  : q <= 23'h232ca6; 
			12'd689  : q <= 23'h000000; 
			12'd690  : q <= 23'h000000; 
			12'd691  : q <= 23'h000000; 
			12'd692  : q <= 23'h000000; 
			12'd693  : q <= 23'h000000; 
			12'd694  : q <= 23'h000000; 
			12'd695  : q <= 23'h000000; 
			12'd696  : q <= 23'h000000; 
			12'd697  : q <= 23'h000000; 
			12'd698  : q <= 23'h000000; 
			12'd699  : q <= 23'h000000; 
			12'd700  : q <= 23'h000000; 
			12'd701  : q <= 23'h000000; 
			12'd702  : q <= 23'h000000; 
			12'd703  : q <= 23'h000000; 
			12'd704  : q <= 23'h000000; 
			12'd705  : q <= 23'h000000; 
			12'd706  : q <= 23'h000000; 
			12'd707  : q <= 23'h000000; 
			12'd708  : q <= 23'h000000; 
			12'd709  : q <= 23'h000000; 
			12'd710  : q <= 23'h23b086; 
			12'd711  : q <= 23'h24b086; 
			12'd712  : q <= 23'h000000; 
			12'd713  : q <= 23'h000000; 
			12'd714  : q <= 23'h000000; 
			12'd715  : q <= 23'h000000; 
			12'd716  : q <= 23'h000000; 
			12'd717  : q <= 23'h000000; 
			12'd718  : q <= 23'h000000; 
			12'd719  : q <= 23'h000000; 
			12'd720  : q <= 23'h000000; 
			12'd721  : q <= 23'h000000; 
			12'd722  : q <= 23'h000000; 
			12'd723  : q <= 23'h000000; 
			12'd724  : q <= 23'h244043; 
			12'd725  : q <= 23'h000000; 
			12'd726  : q <= 23'h000000; 
			12'd727  : q <= 23'h250d41; 
			12'd728  : q <= 23'h000000; 
			12'd729  : q <= 23'h000000; 
			12'd730  : q <= 23'h000000; 
			12'd731  : q <= 23'h000000; 
			12'd732  : q <= 23'h274064; 
			12'd733  : q <= 23'h24c0a3; 
			12'd734  : q <= 23'h000000; 
			12'd735  : q <= 23'h000000; 
			12'd736  : q <= 23'h000000; 
			12'd737  : q <= 23'h000000; 
			12'd738  : q <= 23'h000000; 
			12'd739  : q <= 23'h000000; 
			12'd740  : q <= 23'h000000; 
			12'd741  : q <= 23'h000000; 
			12'd742  : q <= 23'h000000; 
			12'd743  : q <= 23'h000000; 
			12'd744  : q <= 23'h000000; 
			12'd745  : q <= 23'h000000; 
			12'd746  : q <= 23'h000000; 
			12'd747  : q <= 23'h000000; 
			12'd748  : q <= 23'h000000; 
			12'd749  : q <= 23'h21c463; 
			12'd750  : q <= 23'h000000; 
			12'd751  : q <= 23'h000000; 
			12'd752  : q <= 23'h000000; 
			12'd753  : q <= 23'h000000; 
			12'd754  : q <= 23'h000000; 
			12'd755  : q <= 23'h000000; 
			12'd756  : q <= 23'h000000; 
			12'd757  : q <= 23'h000000; 
			12'd758  : q <= 23'h000000; 
			12'd759  : q <= 23'h000000; 
			12'd760  : q <= 23'h000000; 
			12'd761  : q <= 23'h24a8c6; 
			12'd762  : q <= 23'h000000; 
			12'd763  : q <= 23'h000000; 
			12'd764  : q <= 23'h000000; 
			12'd765  : q <= 23'h000000; 
			12'd766  : q <= 23'h000000; 
			12'd767  : q <= 23'h000000; 
			12'd768  : q <= 23'h000000; 
			12'd769  : q <= 23'h000000; 
			12'd770  : q <= 23'h20b523; 
			12'd771  : q <= 23'h000000; 
			12'd772  : q <= 23'h000000; 
			12'd773  : q <= 23'h000000; 
			12'd774  : q <= 23'h000000; 
			12'd775  : q <= 23'h239cc6; 
			12'd776  : q <= 23'h251822; 
			12'd777  : q <= 23'h22a8a1; 
			12'd778  : q <= 23'h000000; 
			12'd779  : q <= 23'h000000; 
			12'd780  : q <= 23'h000000; 
			12'd781  : q <= 23'h000000; 
			12'd782  : q <= 23'h24a462; 
			12'd783  : q <= 23'h000000; 
			12'd784  : q <= 23'h000000; 
			12'd785  : q <= 23'h000000; 
			12'd786  : q <= 23'h000000; 
			12'd787  : q <= 23'h000000; 
			12'd788  : q <= 23'h000000; 
			12'd789  : q <= 23'h000000; 
			12'd790  : q <= 23'h000000; 
			12'd791  : q <= 23'h000000; 
			12'd792  : q <= 23'h000000; 
			12'd793  : q <= 23'h000000; 
			12'd794  : q <= 23'h000000; 
			12'd795  : q <= 23'h234443; 
			12'd796  : q <= 23'h000000; 
			12'd797  : q <= 23'h000000; 
			12'd798  : q <= 23'h271064; 
			12'd799  : q <= 23'h000000; 
			12'd800  : q <= 23'h000000; 
			12'd801  : q <= 23'h251886; 
			12'd802  : q <= 23'h271425; 
			12'd803  : q <= 23'h249883; 
			12'd804  : q <= 23'h271465; 
			12'd805  : q <= 23'h000000; 
			12'd806  : q <= 23'h000000; 
			12'd807  : q <= 23'h000000; 
			12'd808  : q <= 23'h21bce2; 
			12'd809  : q <= 23'h000000; 
			12'd810  : q <= 23'h000000; 
			12'd811  : q <= 23'h000000; 
			12'd812  : q <= 23'h000000; 
			12'd813  : q <= 23'h000000; 
			12'd814  : q <= 23'h2224c5; 
			12'd815  : q <= 23'h000000; 
			12'd816  : q <= 23'h244044; 
			12'd817  : q <= 23'h000000; 
			12'd818  : q <= 23'h000000; 
			12'd819  : q <= 23'h000000; 
			12'd820  : q <= 23'h000000; 
			12'd821  : q <= 23'h000000; 
			12'd822  : q <= 23'h000000; 
			12'd823  : q <= 23'h000000; 
			12'd824  : q <= 23'h000000; 
			12'd825  : q <= 23'h000000; 
			12'd826  : q <= 23'h000000; 
			12'd827  : q <= 23'h000000; 
			12'd828  : q <= 23'h271464; 
			12'd829  : q <= 23'h219464; 
			12'd830  : q <= 23'h209523; 
			12'd831  : q <= 23'h000000; 
			12'd832  : q <= 23'h269443; 
			12'd833  : q <= 23'h000000; 
			12'd834  : q <= 23'h000000; 
			12'd835  : q <= 23'h000000; 
			12'd836  : q <= 23'h269443; 
			12'd837  : q <= 23'h229443; 
			12'd838  : q <= 23'h000000; 
			12'd839  : q <= 23'h000000; 
			12'd840  : q <= 23'h000000; 
			12'd841  : q <= 23'h000000; 
			12'd842  : q <= 23'h000000; 
			12'd843  : q <= 23'h244842; 
			12'd844  : q <= 23'h000000; 
			12'd845  : q <= 23'h000000; 
			12'd846  : q <= 23'h000000; 
			12'd847  : q <= 23'h000000; 
			12'd848  : q <= 23'h000000; 
			12'd849  : q <= 23'h000000; 
			12'd850  : q <= 23'h000000; 
			12'd851  : q <= 23'h000000; 
			12'd852  : q <= 23'h000000; 
			12'd853  : q <= 23'h000000; 
			12'd854  : q <= 23'h000000; 
			12'd855  : q <= 23'h000000; 
			12'd856  : q <= 23'h000000; 
			12'd857  : q <= 23'h000000; 
			12'd858  : q <= 23'h000000; 
			12'd859  : q <= 23'h243021; 
			12'd860  : q <= 23'h000000; 
			12'd861  : q <= 23'h000000; 
			12'd862  : q <= 23'h000000; 
			12'd863  : q <= 23'h000000; 
			12'd864  : q <= 23'h000000; 
			12'd865  : q <= 23'h000000; 
			12'd866  : q <= 23'h000000; 
			12'd867  : q <= 23'h000000; 
			12'd868  : q <= 23'h000000; 
			12'd869  : q <= 23'h000000; 
			12'd870  : q <= 23'h000000; 
			12'd871  : q <= 23'h000000; 
			12'd872  : q <= 23'h000000; 
			12'd873  : q <= 23'h000000; 
			12'd874  : q <= 23'h000000; 
			12'd875  : q <= 23'h000000; 
			12'd876  : q <= 23'h273c45; 
			12'd877  : q <= 23'h000000; 
			12'd878  : q <= 23'h000000; 
			12'd879  : q <= 23'h223c45; 
			12'd880  : q <= 23'h204143; 
			12'd881  : q <= 23'h000000; 
			12'd882  : q <= 23'h20a522; 
			12'd883  : q <= 23'h000000; 
			12'd884  : q <= 23'h212503; 
			12'd885  : q <= 23'h000000; 
			12'd886  : q <= 23'h000000; 
			12'd887  : q <= 23'h248c81; 
			12'd888  : q <= 23'h000000; 
			12'd889  : q <= 23'h000000; 
			12'd890  : q <= 23'h000000; 
			12'd891  : q <= 23'h000000; 
			12'd892  : q <= 23'h000000; 
			12'd893  : q <= 23'h000000; 
			12'd894  : q <= 23'h000000; 
			12'd895  : q <= 23'h000000; 
			12'd896  : q <= 23'h000000; 
			12'd897  : q <= 23'h000000; 
			12'd898  : q <= 23'h000000; 
			12'd899  : q <= 23'h000000; 
			12'd900  : q <= 23'h000000; 
			12'd901  : q <= 23'h000000; 
			12'd902  : q <= 23'h000000; 
			12'd903  : q <= 23'h000000; 
			12'd904  : q <= 23'h000000; 
			12'd905  : q <= 23'h000000; 
			12'd906  : q <= 23'h000000; 
			12'd907  : q <= 23'h000000; 
			12'd908  : q <= 23'h000000; 
			12'd909  : q <= 23'h000000; 
			12'd910  : q <= 23'h000000; 
			12'd911  : q <= 23'h000000; 
			12'd912  : q <= 23'h000000; 
			12'd913  : q <= 23'h000000; 
			12'd914  : q <= 23'h000000; 
			12'd915  : q <= 23'h000000; 
			12'd916  : q <= 23'h000000; 
			12'd917  : q <= 23'h000000; 
			12'd918  : q <= 23'h244862; 
			12'd919  : q <= 23'h000000; 
			12'd920  : q <= 23'h000000; 
			12'd921  : q <= 23'h23ac85; 
			12'd922  : q <= 23'h24ac85; 
			12'd923  : q <= 23'h000000; 
			12'd924  : q <= 23'h000000; 
			12'd925  : q <= 23'h000000; 
			12'd926  : q <= 23'h229425; 
			12'd927  : q <= 23'h000000; 
			12'd928  : q <= 23'h000000; 
			12'd929  : q <= 23'h000000; 
			12'd930  : q <= 23'h000000; 
			12'd931  : q <= 23'h000000; 
			12'd932  : q <= 23'h000000; 
			12'd933  : q <= 23'h000000; 
			12'd934  : q <= 23'h000000; 
			12'd935  : q <= 23'h000000; 
			12'd936  : q <= 23'h000000; 
			12'd937  : q <= 23'h000000; 
			12'd938  : q <= 23'h000000; 
			12'd939  : q <= 23'h000000; 
			12'd940  : q <= 23'h000000; 
			12'd941  : q <= 23'h000000; 
			12'd942  : q <= 23'h000000; 
			12'd943  : q <= 23'h259423; 
			12'd944  : q <= 23'h000000; 
			12'd945  : q <= 23'h000000; 
			12'd946  : q <= 23'h000000; 
			12'd947  : q <= 23'h000000; 
			12'd948  : q <= 23'h000000; 
			12'd949  : q <= 23'h000000; 
			12'd950  : q <= 23'h000000; 
			12'd951  : q <= 23'h000000; 
			12'd952  : q <= 23'h000000; 
			12'd953  : q <= 23'h25bc41; 
			12'd954  : q <= 23'h000000; 
			12'd955  : q <= 23'h000000; 
			12'd956  : q <= 23'h000000; 
			12'd957  : q <= 23'h000000; 
			12'd958  : q <= 23'h000000; 
			12'd959  : q <= 23'h000000; 
			12'd960  : q <= 23'h000000; 
			12'd961  : q <= 23'h000000; 
			12'd962  : q <= 23'h000000; 
			12'd963  : q <= 23'h000000; 
			12'd964  : q <= 23'h000000; 
			12'd965  : q <= 23'h000000; 
			12'd966  : q <= 23'h000000; 
			12'd967  : q <= 23'h000000; 
			12'd968  : q <= 23'h000000; 
			12'd969  : q <= 23'h000000; 
			12'd970  : q <= 23'h000000; 
			12'd971  : q <= 23'h000000; 
			12'd972  : q <= 23'h000000; 
			12'd973  : q <= 23'h000000; 
			12'd974  : q <= 23'h000000; 
			12'd975  : q <= 23'h2294c5; 
			12'd976  : q <= 23'h000000; 
			12'd977  : q <= 23'h000000; 
			12'd978  : q <= 23'h221825; 
			12'd979  : q <= 23'h000000; 
			12'd980  : q <= 23'h000000; 
			12'd981  : q <= 23'h000000; 
			12'd982  : q <= 23'h000000; 
			12'd983  : q <= 23'h213922; 
			12'd984  : q <= 23'h232021; 
			12'd985  : q <= 23'h000000; 
			12'd986  : q <= 23'h20ac29; 
			12'd987  : q <= 23'h209122; 
			12'd988  : q <= 23'h000000; 
			12'd989  : q <= 23'h213922; 
			12'd990  : q <= 23'h24b922; 
			12'd991  : q <= 23'h000000; 
			12'd992  : q <= 23'h000000; 
			12'd993  : q <= 23'h000000; 
			12'd994  : q <= 23'h000000; 
			12'd995  : q <= 23'h000000; 
			12'd996  : q <= 23'h000000; 
			12'd997  : q <= 23'h259024; 
			12'd998  : q <= 23'h21b866; 
			12'd999  : q <= 23'h000000; 
			12'd1000 : q <= 23'h000000; 
			12'd1001 : q <= 23'h000000; 
			12'd1002 : q <= 23'h000000; 
			12'd1003 : q <= 23'h000000; 
			12'd1004 : q <= 23'h251444; 
			12'd1005 : q <= 23'h000000; 
			12'd1006 : q <= 23'h000000; 
			12'd1007 : q <= 23'h000000; 
			12'd1008 : q <= 23'h000000; 
			12'd1009 : q <= 23'h000000; 
			12'd1010 : q <= 23'h000000; 
			12'd1011 : q <= 23'h000000; 
			12'd1012 : q <= 23'h000000; 
			12'd1013 : q <= 23'h20a525; 
			12'd1014 : q <= 23'h000000; 
			12'd1015 : q <= 23'h000000; 
			12'd1016 : q <= 23'h000000; 
			12'd1017 : q <= 23'h000000; 
			12'd1018 : q <= 23'h000000; 
			12'd1019 : q <= 23'h000000; 
			12'd1020 : q <= 23'h000000; 
			12'd1021 : q <= 23'h000000; 
			12'd1022 : q <= 23'h000000; 
			12'd1023 : q <= 23'h291c24; 
			12'd1024 : q <= 23'h209c24; 
			12'd1025 : q <= 23'h21b0e5; 
			12'd1026 : q <= 23'h000000; 
			12'd1027 : q <= 23'h000000; 
			12'd1028 : q <= 23'h000000; 
			12'd1029 : q <= 23'h000000; 
			12'd1030 : q <= 23'h000000; 
			12'd1031 : q <= 23'h000000; 
			12'd1032 : q <= 23'h000000; 
			12'd1033 : q <= 23'h000000; 
			12'd1034 : q <= 23'h000000; 
			12'd1035 : q <= 23'h000000; 
			12'd1036 : q <= 23'h219465; 
			12'd1037 : q <= 23'h000000; 
			12'd1038 : q <= 23'h000000; 
			12'd1039 : q <= 23'h000000; 
			12'd1040 : q <= 23'h000000; 
			12'd1041 : q <= 23'h2330e1; 
			12'd1042 : q <= 23'h249821; 
			12'd1043 : q <= 23'h000000; 
			12'd1044 : q <= 23'h000000; 
			12'd1045 : q <= 23'h000000; 
			12'd1046 : q <= 23'h000000; 
			12'd1047 : q <= 23'h000000; 
			12'd1048 : q <= 23'h000000; 
			12'd1049 : q <= 23'h244043; 
			12'd1050 : q <= 23'h000000; 
			12'd1051 : q <= 23'h000000; 
			12'd1052 : q <= 23'h231023; 
			12'd1053 : q <= 23'h000000; 
			12'd1054 : q <= 23'h000000; 
			12'd1055 : q <= 23'h000000; 
			12'd1056 : q <= 23'h000000; 
			12'd1057 : q <= 23'h2424e5; 
			12'd1058 : q <= 23'h25b467; 
			12'd1059 : q <= 23'h233467; 
			12'd1060 : q <= 23'h000000; 
			12'd1061 : q <= 23'h000000; 
			12'd1062 : q <= 23'h2314e2; 
			12'd1063 : q <= 23'h000000; 
			12'd1064 : q <= 23'h000000; 
			12'd1065 : q <= 23'h000000; 
			12'd1066 : q <= 23'h000000; 
			12'd1067 : q <= 23'h242462; 
			12'd1068 : q <= 23'h000000; 
			12'd1069 : q <= 23'h000000; 
			12'd1070 : q <= 23'h000000; 
			12'd1071 : q <= 23'h000000; 
			12'd1072 : q <= 23'h000000; 
			12'd1073 : q <= 23'h000000; 
			12'd1074 : q <= 23'h000000; 
			12'd1075 : q <= 23'h000000; 
			12'd1076 : q <= 23'h000000; 
			12'd1077 : q <= 23'h000000; 
			12'd1078 : q <= 23'h000000; 
			12'd1079 : q <= 23'h000000; 
			12'd1080 : q <= 23'h000000; 
			12'd1081 : q <= 23'h000000; 
			12'd1082 : q <= 23'h000000; 
			12'd1083 : q <= 23'h000000; 
			12'd1084 : q <= 23'h000000; 
			12'd1085 : q <= 23'h000000; 
			12'd1086 : q <= 23'h000000; 
			12'd1087 : q <= 23'h000000; 
			12'd1088 : q <= 23'h251c41; 
			12'd1089 : q <= 23'h241c41; 
			12'd1090 : q <= 23'h000000; 
			12'd1091 : q <= 23'h000000; 
			12'd1092 : q <= 23'h000000; 
			12'd1093 : q <= 23'h000000; 
			12'd1094 : q <= 23'h211522; 
			12'd1095 : q <= 23'h000000; 
			12'd1096 : q <= 23'h000000; 
			12'd1097 : q <= 23'h000000; 
			12'd1098 : q <= 23'h000000; 
			12'd1099 : q <= 23'h000000; 
			12'd1100 : q <= 23'h000000; 
			12'd1101 : q <= 23'h000000; 
			12'd1102 : q <= 23'h000000; 
			12'd1103 : q <= 23'h000000; 
			12'd1104 : q <= 23'h000000; 
			12'd1105 : q <= 23'h000000; 
			12'd1106 : q <= 23'h000000; 
			12'd1107 : q <= 23'h000000; 
			12'd1108 : q <= 23'h000000; 
			12'd1109 : q <= 23'h253483; 
			12'd1110 : q <= 23'h000000; 
			12'd1111 : q <= 23'h000000; 
			12'd1112 : q <= 23'h000000; 
			12'd1113 : q <= 23'h000000; 
			12'd1114 : q <= 23'h000000; 
			12'd1115 : q <= 23'h000000; 
			12'd1116 : q <= 23'h000000; 
			12'd1117 : q <= 23'h000000; 
			12'd1118 : q <= 23'h000000; 
			12'd1119 : q <= 23'h000000; 
			12'd1120 : q <= 23'h000000; 
			12'd1121 : q <= 23'h000000; 
			12'd1122 : q <= 23'h20cd21; 
			12'd1123 : q <= 23'h000000; 
			12'd1124 : q <= 23'h000000; 
			12'd1125 : q <= 23'h000000; 
			12'd1126 : q <= 23'h000000; 
			12'd1127 : q <= 23'h000000; 
			12'd1128 : q <= 23'h000000; 
			12'd1129 : q <= 23'h000000; 
			12'd1130 : q <= 23'h000000; 
			12'd1131 : q <= 23'h000000; 
			12'd1132 : q <= 23'h000000; 
			12'd1133 : q <= 23'h000000; 
			12'd1134 : q <= 23'h000000; 
			12'd1135 : q <= 23'h000000; 
			12'd1136 : q <= 23'h000000; 
			12'd1137 : q <= 23'h000000; 
			12'd1138 : q <= 23'h000000; 
			12'd1139 : q <= 23'h000000; 
			12'd1140 : q <= 23'h261481; 
			12'd1141 : q <= 23'h221481; 
			12'd1142 : q <= 23'h000000; 
			12'd1143 : q <= 23'h000000; 
			12'd1144 : q <= 23'h000000; 
			12'd1145 : q <= 23'h000000; 
			12'd1146 : q <= 23'h262044; 
			12'd1147 : q <= 23'h23a021; 
			12'd1148 : q <= 23'h000000; 
			12'd1149 : q <= 23'h000000; 
			12'd1150 : q <= 23'h000000; 
			12'd1151 : q <= 23'h000000; 
			12'd1152 : q <= 23'h000000; 
			12'd1153 : q <= 23'h000000; 
			12'd1154 : q <= 23'h000000; 
			12'd1155 : q <= 23'h000000; 
			12'd1156 : q <= 23'h000000; 
			12'd1157 : q <= 23'h000000; 
			12'd1158 : q <= 23'h000000; 
			12'd1159 : q <= 23'h000000; 
			12'd1160 : q <= 23'h213102; 
			12'd1161 : q <= 23'h000000; 
			12'd1162 : q <= 23'h000000; 
			12'd1163 : q <= 23'h000000; 
			12'd1164 : q <= 23'h000000; 
			12'd1165 : q <= 23'h251886; 
			12'd1166 : q <= 23'h26a021; 
			12'd1167 : q <= 23'h000000; 
			12'd1168 : q <= 23'h000000; 
			12'd1169 : q <= 23'h000000; 
			12'd1170 : q <= 23'h000000; 
			12'd1171 : q <= 23'h000000; 
			12'd1172 : q <= 23'h000000; 
			12'd1173 : q <= 23'h000000; 
			12'd1174 : q <= 23'h000000; 
			12'd1175 : q <= 23'h000000; 
			12'd1176 : q <= 23'h000000; 
			12'd1177 : q <= 23'h000000; 
			12'd1178 : q <= 23'h202543; 
			12'd1179 : q <= 23'h221c21; 
			12'd1180 : q <= 23'h279c21; 
			12'd1181 : q <= 23'h221c21; 
			12'd1182 : q <= 23'h000000; 
			12'd1183 : q <= 23'h252905; 
			12'd1184 : q <= 23'h000000; 
			12'd1185 : q <= 23'h000000; 
			12'd1186 : q <= 23'h000000; 
			12'd1187 : q <= 23'h000000; 
			12'd1188 : q <= 23'h000000; 
			12'd1189 : q <= 23'h000000; 
			12'd1190 : q <= 23'h000000; 
			12'd1191 : q <= 23'h000000; 
			12'd1192 : q <= 23'h000000; 
			12'd1193 : q <= 23'h000000; 
			12'd1194 : q <= 23'h26a462; 
			12'd1195 : q <= 23'h000000; 
			12'd1196 : q <= 23'h000000; 
			12'd1197 : q <= 23'h241463; 
			12'd1198 : q <= 23'h24c862; 
			12'd1199 : q <= 23'h000000; 
			12'd1200 : q <= 23'h000000; 
			12'd1201 : q <= 23'h000000; 
			12'd1202 : q <= 23'h000000; 
			12'd1203 : q <= 23'h000000; 
			12'd1204 : q <= 23'h23b863; 
			12'd1205 : q <= 23'h000000; 
			12'd1206 : q <= 23'h000000; 
			12'd1207 : q <= 23'h000000; 
			12'd1208 : q <= 23'h000000; 
			12'd1209 : q <= 23'h000000; 
			12'd1210 : q <= 23'h000000; 
			12'd1211 : q <= 23'h000000; 
			12'd1212 : q <= 23'h000000; 
			12'd1213 : q <= 23'h000000; 
			12'd1214 : q <= 23'h000000; 
			12'd1215 : q <= 23'h000000; 
			12'd1216 : q <= 23'h000000; 
			12'd1217 : q <= 23'h000000; 
			12'd1218 : q <= 23'h000000; 
			12'd1219 : q <= 23'h000000; 
			12'd1220 : q <= 23'h000000; 
			12'd1221 : q <= 23'h000000; 
			12'd1222 : q <= 23'h000000; 
			12'd1223 : q <= 23'h000000; 
			12'd1224 : q <= 23'h000000; 
			12'd1225 : q <= 23'h000000; 
			12'd1226 : q <= 23'h000000; 
			12'd1227 : q <= 23'h000000; 
			12'd1228 : q <= 23'h000000; 
			12'd1229 : q <= 23'h000000; 
			12'd1230 : q <= 23'h000000; 
			12'd1231 : q <= 23'h000000; 
			12'd1232 : q <= 23'h000000; 
			12'd1233 : q <= 23'h251886; 
			12'd1234 : q <= 23'h000000; 
			12'd1235 : q <= 23'h000000; 
			12'd1236 : q <= 23'h000000; 
			12'd1237 : q <= 23'h000000; 
			12'd1238 : q <= 23'h24b461; 
			12'd1239 : q <= 23'h000000; 
			12'd1240 : q <= 23'h259c21; 
			12'd1241 : q <= 23'h000000; 
			12'd1242 : q <= 23'h259c21; 
			12'd1243 : q <= 23'h000000; 
			12'd1244 : q <= 23'h000000; 
			12'd1245 : q <= 23'h000000; 
			12'd1246 : q <= 23'h000000; 
			12'd1247 : q <= 23'h000000; 
			12'd1248 : q <= 23'h000000; 
			12'd1249 : q <= 23'h000000; 
			12'd1250 : q <= 23'h000000; 
			12'd1251 : q <= 23'h000000; 
			12'd1252 : q <= 23'h000000; 
			12'd1253 : q <= 23'h000000; 
			12'd1254 : q <= 23'h264021; 
			12'd1255 : q <= 23'h000000; 
			12'd1256 : q <= 23'h000000; 
			12'd1257 : q <= 23'h000000; 
			12'd1258 : q <= 23'h000000; 
			12'd1259 : q <= 23'h000000; 
			12'd1260 : q <= 23'h000000; 
			12'd1261 : q <= 23'h229c26; 
			12'd1262 : q <= 23'h25c463; 
			12'd1263 : q <= 23'h234463; 
			12'd1264 : q <= 23'h000000; 
			12'd1265 : q <= 23'h000000; 
			12'd1266 : q <= 23'h000000; 
			12'd1267 : q <= 23'h000000; 
			12'd1268 : q <= 23'h000000; 
			12'd1269 : q <= 23'h23c021; 
			12'd1270 : q <= 23'h233883; 
			12'd1271 : q <= 23'h241c21; 
			12'd1272 : q <= 23'h211503; 
			12'd1273 : q <= 23'h000000; 
			12'd1274 : q <= 23'h000000; 
			12'd1275 : q <= 23'h000000; 
			12'd1276 : q <= 23'h000000; 
			12'd1277 : q <= 23'h000000; 
			12'd1278 : q <= 23'h000000; 
			12'd1279 : q <= 23'h21ac49; 
			12'd1280 : q <= 23'h000000; 
			12'd1281 : q <= 23'h000000; 
			12'd1282 : q <= 23'h000000; 
			12'd1283 : q <= 23'h000000; 
			12'd1284 : q <= 23'h000000; 
			12'd1285 : q <= 23'h000000; 
			12'd1286 : q <= 23'h000000; 
			12'd1287 : q <= 23'h000000; 
			12'd1288 : q <= 23'h262883; 
			12'd1289 : q <= 23'h222883; 
			12'd1290 : q <= 23'h291c25; 
			12'd1291 : q <= 23'h000000; 
			12'd1292 : q <= 23'h000000; 
			12'd1293 : q <= 23'h244021; 
			12'd1294 : q <= 23'h000000; 
			12'd1295 : q <= 23'h000000; 
			12'd1296 : q <= 23'h000000; 
			12'd1297 : q <= 23'h000000; 
			12'd1298 : q <= 23'h000000; 
			12'd1299 : q <= 23'h000000; 
			12'd1300 : q <= 23'h000000; 
			12'd1301 : q <= 23'h000000; 
			12'd1302 : q <= 23'h000000; 
			12'd1303 : q <= 23'h243821; 
			12'd1304 : q <= 23'h2234e2; 
			12'd1305 : q <= 23'h000000; 
			12'd1306 : q <= 23'h25cc21; 
			12'd1307 : q <= 23'h244c21; 
			12'd1308 : q <= 23'h000000; 
			12'd1309 : q <= 23'h000000; 
			12'd1310 : q <= 23'h244044; 
			12'd1311 : q <= 23'h000000; 
			12'd1312 : q <= 23'h000000; 
			12'd1313 : q <= 23'h000000; 
			12'd1314 : q <= 23'h000000; 
			12'd1315 : q <= 23'h000000; 
			12'd1316 : q <= 23'h000000; 
			12'd1317 : q <= 23'h000000; 
			12'd1318 : q <= 23'h000000; 
			12'd1319 : q <= 23'h000000; 
			12'd1320 : q <= 23'h25b021; 
			12'd1321 : q <= 23'h000000; 
			12'd1322 : q <= 23'h25b021; 
			12'd1323 : q <= 23'h000000; 
			12'd1324 : q <= 23'h25b021; 
			12'd1325 : q <= 23'h000000; 
			12'd1326 : q <= 23'h25b021; 
			12'd1327 : q <= 23'h243021; 
			12'd1328 : q <= 23'h000000; 
			12'd1329 : q <= 23'h000000; 
			12'd1330 : q <= 23'h000000; 
			12'd1331 : q <= 23'h000000; 
			12'd1332 : q <= 23'h000000; 
			12'd1333 : q <= 23'h000000; 
			12'd1334 : q <= 23'h000000; 
			12'd1335 : q <= 23'h254024; 
			12'd1336 : q <= 23'h25a021; 
			12'd1337 : q <= 23'h000000; 
			12'd1338 : q <= 23'h000000; 
			12'd1339 : q <= 23'h000000; 
			12'd1340 : q <= 23'h000000; 
			12'd1341 : q <= 23'h000000; 
			12'd1342 : q <= 23'h000000; 
			12'd1343 : q <= 23'h000000; 
			12'd1344 : q <= 23'h000000; 
			12'd1345 : q <= 23'h000000; 
			12'd1346 : q <= 23'h000000; 
			12'd1347 : q <= 23'h000000; 
			12'd1348 : q <= 23'h263421; 
			12'd1349 : q <= 23'h23b421; 
			12'd1350 : q <= 23'h242841; 
			12'd1351 : q <= 23'h221c21; 
			12'd1352 : q <= 23'h000000; 
			12'd1353 : q <= 23'h000000; 
			12'd1354 : q <= 23'h000000; 
			12'd1355 : q <= 23'h000000; 
			12'd1356 : q <= 23'h000000; 
			12'd1357 : q <= 23'h222462; 
			12'd1358 : q <= 23'h000000; 
			12'd1359 : q <= 23'h000000; 
			12'd1360 : q <= 23'h000000; 
			12'd1361 : q <= 23'h000000; 
			12'd1362 : q <= 23'h000000; 
			12'd1363 : q <= 23'h000000; 
			12'd1364 : q <= 23'h000000; 
			12'd1365 : q <= 23'h000000; 
			12'd1366 : q <= 23'h000000; 
			12'd1367 : q <= 23'h000000; 
			12'd1368 : q <= 23'h000000; 
			12'd1369 : q <= 23'h000000; 
			12'd1370 : q <= 23'h000000; 
			12'd1371 : q <= 23'h000000; 
			12'd1372 : q <= 23'h000000; 
			12'd1373 : q <= 23'h000000; 
			12'd1374 : q <= 23'h000000; 
			12'd1375 : q <= 23'h000000; 
			12'd1376 : q <= 23'h000000; 
			12'd1377 : q <= 23'h000000; 
			12'd1378 : q <= 23'h000000; 
			12'd1379 : q <= 23'h000000; 
			12'd1380 : q <= 23'h000000; 
			12'd1381 : q <= 23'h000000; 
			12'd1382 : q <= 23'h000000; 
			12'd1383 : q <= 23'h000000; 
			12'd1384 : q <= 23'h000000; 
			12'd1385 : q <= 23'h000000; 
			12'd1386 : q <= 23'h000000; 
			12'd1387 : q <= 23'h000000; 
			12'd1388 : q <= 23'h250c43; 
			12'd1389 : q <= 23'h000000; 
			12'd1390 : q <= 23'h260481; 
			12'd1391 : q <= 23'h000000; 
			12'd1392 : q <= 23'h28b025; 
			12'd1393 : q <= 23'h213025; 
			12'd1394 : q <= 23'h000000; 
			12'd1395 : q <= 23'h000000; 
			12'd1396 : q <= 23'h000000; 
			12'd1397 : q <= 23'h220481; 
			12'd1398 : q <= 23'h000000; 
			12'd1399 : q <= 23'h000000; 
			12'd1400 : q <= 23'h000000; 
			12'd1401 : q <= 23'h000000; 
			12'd1402 : q <= 23'h000000; 
			12'd1403 : q <= 23'h000000; 
			12'd1404 : q <= 23'h000000; 
			12'd1405 : q <= 23'h000000; 
			12'd1406 : q <= 23'h000000; 
			12'd1407 : q <= 23'h000000; 
			12'd1408 : q <= 23'h000000; 
			12'd1409 : q <= 23'h000000; 
			12'd1410 : q <= 23'h000000; 
			12'd1411 : q <= 23'h000000; 
			12'd1412 : q <= 23'h000000; 
			12'd1413 : q <= 23'h000000; 
			12'd1414 : q <= 23'h201543; 
			12'd1415 : q <= 23'h000000; 
			12'd1416 : q <= 23'h000000; 
			12'd1417 : q <= 23'h000000; 
			12'd1418 : q <= 23'h000000; 
			12'd1419 : q <= 23'h000000; 
			12'd1420 : q <= 23'h283c45; 
			12'd1421 : q <= 23'h000000; 
			12'd1422 : q <= 23'h000000; 
			12'd1423 : q <= 23'h213c45; 
			12'd1424 : q <= 23'h000000; 
			12'd1425 : q <= 23'h000000; 
			12'd1426 : q <= 23'h000000; 
			12'd1427 : q <= 23'h000000; 
			12'd1428 : q <= 23'h000000; 
			12'd1429 : q <= 23'h000000; 
			12'd1430 : q <= 23'h000000; 
			12'd1431 : q <= 23'h000000; 
			12'd1432 : q <= 23'h000000; 
			12'd1433 : q <= 23'h000000; 
			12'd1434 : q <= 23'h000000; 
			12'd1435 : q <= 23'h000000; 
			12'd1436 : q <= 23'h000000; 
			12'd1437 : q <= 23'h000000; 
			12'd1438 : q <= 23'h000000; 
			12'd1439 : q <= 23'h000000; 
			12'd1440 : q <= 23'h000000; 
			12'd1441 : q <= 23'h000000; 
			12'd1442 : q <= 23'h000000; 
			12'd1443 : q <= 23'h000000; 
			12'd1444 : q <= 23'h000000; 
			12'd1445 : q <= 23'h000000; 
			12'd1446 : q <= 23'h000000; 
			12'd1447 : q <= 23'h000000; 
			12'd1448 : q <= 23'h000000; 
			12'd1449 : q <= 23'h000000; 
			12'd1450 : q <= 23'h258c23; 
			12'd1451 : q <= 23'h240c23; 
			12'd1452 : q <= 23'h000000; 
			12'd1453 : q <= 23'h000000; 
			12'd1454 : q <= 23'h000000; 
			12'd1455 : q <= 23'h000000; 
			12'd1456 : q <= 23'h211104; 
			12'd1457 : q <= 23'h000000; 
			12'd1458 : q <= 23'h000000; 
			12'd1459 : q <= 23'h000000; 
			12'd1460 : q <= 23'h000000; 
			12'd1461 : q <= 23'h000000; 
			12'd1462 : q <= 23'h000000; 
			12'd1463 : q <= 23'h24a502; 
			12'd1464 : q <= 23'h000000; 
			12'd1465 : q <= 23'h000000; 
			12'd1466 : q <= 23'h2228e5; 
			12'd1467 : q <= 23'h000000; 
			12'd1468 : q <= 23'h000000; 
			12'd1469 : q <= 23'h000000; 
			12'd1470 : q <= 23'h000000; 
			12'd1471 : q <= 23'h000000; 
			12'd1472 : q <= 23'h000000; 
			12'd1473 : q <= 23'h000000; 
			12'd1474 : q <= 23'h000000; 
			12'd1475 : q <= 23'h000000; 
			12'd1476 : q <= 23'h000000; 
			12'd1477 : q <= 23'h000000; 
			12'd1478 : q <= 23'h000000; 
			12'd1479 : q <= 23'h000000; 
			12'd1480 : q <= 23'h000000; 
			12'd1481 : q <= 23'h000000; 
			12'd1482 : q <= 23'h000000; 
			12'd1483 : q <= 23'h000000; 
			12'd1484 : q <= 23'h000000; 
			12'd1485 : q <= 23'h000000; 
			12'd1486 : q <= 23'h000000; 
			12'd1487 : q <= 23'h000000; 
			12'd1488 : q <= 23'h000000; 
			12'd1489 : q <= 23'h000000; 
			12'd1490 : q <= 23'h000000; 
			12'd1491 : q <= 23'h000000; 
			12'd1492 : q <= 23'h24cc81; 
			12'd1493 : q <= 23'h000000; 
			12'd1494 : q <= 23'h000000; 
			12'd1495 : q <= 23'h000000; 
			12'd1496 : q <= 23'h000000; 
			12'd1497 : q <= 23'h000000; 
			12'd1498 : q <= 23'h2214e4; 
			12'd1499 : q <= 23'h223048; 
			12'd1500 : q <= 23'h000000; 
			12'd1501 : q <= 23'h24aca6; 
			12'd1502 : q <= 23'h000000; 
			12'd1503 : q <= 23'h000000; 
			12'd1504 : q <= 23'h261c45; 
			12'd1505 : q <= 23'h000000; 
			12'd1506 : q <= 23'h210521; 
			12'd1507 : q <= 23'h248521; 
			12'd1508 : q <= 23'h26c043; 
			12'd1509 : q <= 23'h22c043; 
			12'd1510 : q <= 23'h000000; 
			12'd1511 : q <= 23'h2538a5; 
			12'd1512 : q <= 23'h259441; 
			12'd1513 : q <= 23'h000000; 
			12'd1514 : q <= 23'h261c45; 
			12'd1515 : q <= 23'h000000; 
			12'd1516 : q <= 23'h000000; 
			12'd1517 : q <= 23'h000000; 
			12'd1518 : q <= 23'h261c45; 
			12'd1519 : q <= 23'h231c45; 
			12'd1520 : q <= 23'h259441; 
			12'd1521 : q <= 23'h000000; 
			12'd1522 : q <= 23'h259441; 
			12'd1523 : q <= 23'h000000; 
			12'd1524 : q <= 23'h259441; 
			12'd1525 : q <= 23'h239441; 
			12'd1526 : q <= 23'h269826; 
			12'd1527 : q <= 23'h000000; 
			12'd1528 : q <= 23'h000000; 
			12'd1529 : q <= 23'h000000; 
			12'd1530 : q <= 23'h000000; 
			12'd1531 : q <= 23'h000000; 
			12'd1532 : q <= 23'h242462; 
			12'd1533 : q <= 23'h000000; 
			12'd1534 : q <= 23'h000000; 
			12'd1535 : q <= 23'h000000; 
			12'd1536 : q <= 23'h231c45; 
			12'd1537 : q <= 23'h000000; 
			12'd1538 : q <= 23'h000000; 
			12'd1539 : q <= 23'h000000; 
			12'd1540 : q <= 23'h000000; 
			12'd1541 : q <= 23'h000000; 
			12'd1542 : q <= 23'h000000; 
			12'd1543 : q <= 23'h000000; 
			12'd1544 : q <= 23'h000000; 
			12'd1545 : q <= 23'h000000; 
			12'd1546 : q <= 23'h000000; 
			12'd1547 : q <= 23'h000000; 
			12'd1548 : q <= 23'h000000; 
			12'd1549 : q <= 23'h000000; 
			12'd1550 : q <= 23'h221485; 
			12'd1551 : q <= 23'h000000; 
			12'd1552 : q <= 23'h000000; 
			12'd1553 : q <= 23'h000000; 
			12'd1554 : q <= 23'h000000; 
			12'd1555 : q <= 23'h000000; 
			12'd1556 : q <= 23'h000000; 
			12'd1557 : q <= 23'h000000; 
			12'd1558 : q <= 23'h000000; 
			12'd1559 : q <= 23'h000000; 
			12'd1560 : q <= 23'h000000; 
			12'd1561 : q <= 23'h000000; 
			12'd1562 : q <= 23'h000000; 
			12'd1563 : q <= 23'h000000; 
			12'd1564 : q <= 23'h000000; 
			12'd1565 : q <= 23'h000000; 
			12'd1566 : q <= 23'h000000; 
			12'd1567 : q <= 23'h000000; 
			12'd1568 : q <= 23'h000000; 
			12'd1569 : q <= 23'h000000; 
			12'd1570 : q <= 23'h000000; 
			12'd1571 : q <= 23'h000000; 
			12'd1572 : q <= 23'h000000; 
			12'd1573 : q <= 23'h000000; 
			12'd1574 : q <= 23'h000000; 
			12'd1575 : q <= 23'h000000; 
			12'd1576 : q <= 23'h000000; 
			12'd1577 : q <= 23'h000000; 
			12'd1578 : q <= 23'h000000; 
			12'd1579 : q <= 23'h000000; 
			12'd1580 : q <= 23'h000000; 
			12'd1581 : q <= 23'h000000; 
			12'd1582 : q <= 23'h000000; 
			12'd1583 : q <= 23'h000000; 
			12'd1584 : q <= 23'h000000; 
			12'd1585 : q <= 23'h000000; 
			12'd1586 : q <= 23'h000000; 
			12'd1587 : q <= 23'h000000; 
			12'd1588 : q <= 23'h000000; 
			12'd1589 : q <= 23'h000000; 
			12'd1590 : q <= 23'h000000; 
			12'd1591 : q <= 23'h000000; 
			12'd1592 : q <= 23'h252cc6; 
			12'd1593 : q <= 23'h233484; 
			12'd1594 : q <= 23'h000000; 
			12'd1595 : q <= 23'h000000; 
			12'd1596 : q <= 23'h000000; 
			12'd1597 : q <= 23'h000000; 
			12'd1598 : q <= 23'h000000; 
			12'd1599 : q <= 23'h000000; 
			12'd1600 : q <= 23'h24b842; 
			12'd1601 : q <= 23'h253021; 
			12'd1602 : q <= 23'h000000; 
			12'd1603 : q <= 23'h253021; 
			12'd1604 : q <= 23'h000000; 
			12'd1605 : q <= 23'h253021; 
			12'd1606 : q <= 23'h24b021; 
			12'd1607 : q <= 23'h000000; 
			12'd1608 : q <= 23'h000000; 
			12'd1609 : q <= 23'h000000; 
			12'd1610 : q <= 23'h000000; 
			12'd1611 : q <= 23'h250441; 
			12'd1612 : q <= 23'h000000; 
			12'd1613 : q <= 23'h243c44; 
			12'd1614 : q <= 23'h000000; 
			12'd1615 : q <= 23'h000000; 
			12'd1616 : q <= 23'h21b026; 
			12'd1617 : q <= 23'h000000; 
			12'd1618 : q <= 23'h000000; 
			12'd1619 : q <= 23'h000000; 
			12'd1620 : q <= 23'h000000; 
			12'd1621 : q <= 23'h248c41; 
			12'd1622 : q <= 23'h000000; 
			12'd1623 : q <= 23'h000000; 
			12'd1624 : q <= 23'h000000; 
			12'd1625 : q <= 23'h000000; 
			12'd1626 : q <= 23'h000000; 
			12'd1627 : q <= 23'h000000; 
			12'd1628 : q <= 23'h000000; 
			12'd1629 : q <= 23'h000000; 
			12'd1630 : q <= 23'h000000; 
			12'd1631 : q <= 23'h000000; 
			12'd1632 : q <= 23'h000000; 
			12'd1633 : q <= 23'h248861; 
			12'd1634 : q <= 23'h000000; 
			12'd1635 : q <= 23'h243441; 
			12'd1636 : q <= 23'h2328a1; 
			12'd1637 : q <= 23'h000000; 
			12'd1638 : q <= 23'h000000; 
			12'd1639 : q <= 23'h000000; 
			12'd1640 : q <= 23'h000000; 
			12'd1641 : q <= 23'h000000; 
			12'd1642 : q <= 23'h24a081; 
			12'd1643 : q <= 23'h000000; 
			12'd1644 : q <= 23'h000000; 
			12'd1645 : q <= 23'h000000; 
			12'd1646 : q <= 23'h000000; 
			12'd1647 : q <= 23'h000000; 
			12'd1648 : q <= 23'h000000; 
			12'd1649 : q <= 23'h000000; 
			12'd1650 : q <= 23'h000000; 
			12'd1651 : q <= 23'h000000; 
			12'd1652 : q <= 23'h000000; 
			12'd1653 : q <= 23'h000000; 
			12'd1654 : q <= 23'h000000; 
			12'd1655 : q <= 23'h24a464; 
			12'd1656 : q <= 23'h242464; 
			12'd1657 : q <= 23'h000000; 
			12'd1658 : q <= 23'h000000; 
			12'd1659 : q <= 23'h000000; 
			12'd1660 : q <= 23'h000000; 
			12'd1661 : q <= 23'h000000; 
			12'd1662 : q <= 23'h000000; 
			12'd1663 : q <= 23'h000000; 
			12'd1664 : q <= 23'h000000; 
			12'd1665 : q <= 23'h000000; 
			12'd1666 : q <= 23'h000000; 
			12'd1667 : q <= 23'h000000; 
			12'd1668 : q <= 23'h000000; 
			12'd1669 : q <= 23'h000000; 
			12'd1670 : q <= 23'h000000; 
			12'd1671 : q <= 23'h000000; 
			12'd1672 : q <= 23'h000000; 
			12'd1673 : q <= 23'h26b465; 
			12'd1674 : q <= 23'h000000; 
			12'd1675 : q <= 23'h263021; 
			12'd1676 : q <= 23'h000000; 
			12'd1677 : q <= 23'h000000; 
			12'd1678 : q <= 23'h000000; 
			12'd1679 : q <= 23'h000000; 
			12'd1680 : q <= 23'h000000; 
			12'd1681 : q <= 23'h000000; 
			12'd1682 : q <= 23'h23b021; 
			12'd1683 : q <= 23'h000000; 
			12'd1684 : q <= 23'h000000; 
			12'd1685 : q <= 23'h274064; 
			12'd1686 : q <= 23'h000000; 
			12'd1687 : q <= 23'h000000; 
			12'd1688 : q <= 23'h000000; 
			12'd1689 : q <= 23'h000000; 
			12'd1690 : q <= 23'h000000; 
			12'd1691 : q <= 23'h222cc2; 
			12'd1692 : q <= 23'h244061; 
			12'd1693 : q <= 23'h000000; 
			12'd1694 : q <= 23'h253941; 
			12'd1695 : q <= 23'h2234c4; 
			12'd1696 : q <= 23'h000000; 
			12'd1697 : q <= 23'h000000; 
			12'd1698 : q <= 23'h253421; 
			12'd1699 : q <= 23'h2234e2; 
			12'd1700 : q <= 23'h000000; 
			12'd1701 : q <= 23'h000000; 
			12'd1702 : q <= 23'h000000; 
			12'd1703 : q <= 23'h26b866; 
			12'd1704 : q <= 23'h223866; 
			12'd1705 : q <= 23'h000000; 
			12'd1706 : q <= 23'h24b482; 
			12'd1707 : q <= 23'h254882; 
			12'd1708 : q <= 23'h000000; 
			12'd1709 : q <= 23'h000000; 
			12'd1710 : q <= 23'h000000; 
			12'd1711 : q <= 23'h000000; 
			12'd1712 : q <= 23'h000000; 
			12'd1713 : q <= 23'h000000; 
			12'd1714 : q <= 23'h000000; 
			12'd1715 : q <= 23'h000000; 
			12'd1716 : q <= 23'h000000; 
			12'd1717 : q <= 23'h000000; 
			12'd1718 : q <= 23'h000000; 
			12'd1719 : q <= 23'h2444a2; 
			12'd1720 : q <= 23'h000000; 
			12'd1721 : q <= 23'h000000; 
			12'd1722 : q <= 23'h000000; 
			12'd1723 : q <= 23'h000000; 
			12'd1724 : q <= 23'h000000; 
			12'd1725 : q <= 23'h000000; 
			12'd1726 : q <= 23'h000000; 
			12'd1727 : q <= 23'h000000; 
			12'd1728 : q <= 23'h000000; 
			12'd1729 : q <= 23'h000000; 
			12'd1730 : q <= 23'h000000; 
			12'd1731 : q <= 23'h000000; 
			12'd1732 : q <= 23'h000000; 
			12'd1733 : q <= 23'h000000; 
			12'd1734 : q <= 23'h000000; 
			12'd1735 : q <= 23'h000000; 
			12'd1736 : q <= 23'h000000; 
			12'd1737 : q <= 23'h000000; 
			12'd1738 : q <= 23'h000000; 
			12'd1739 : q <= 23'h000000; 
			12'd1740 : q <= 23'h000000; 
			12'd1741 : q <= 23'h2314c3; 
			12'd1742 : q <= 23'h000000; 
			12'd1743 : q <= 23'h2214e3; 
			12'd1744 : q <= 23'h000000; 
			12'd1745 : q <= 23'h000000; 
			12'd1746 : q <= 23'h000000; 
			12'd1747 : q <= 23'h000000; 
			12'd1748 : q <= 23'h000000; 
			12'd1749 : q <= 23'h000000; 
			12'd1750 : q <= 23'h000000; 
			12'd1751 : q <= 23'h000000; 
			12'd1752 : q <= 23'h000000; 
			12'd1753 : q <= 23'h000000; 
			12'd1754 : q <= 23'h000000; 
			12'd1755 : q <= 23'h000000; 
			12'd1756 : q <= 23'h000000; 
			12'd1757 : q <= 23'h000000; 
			12'd1758 : q <= 23'h000000; 
			12'd1759 : q <= 23'h000000; 
			12'd1760 : q <= 23'h000000; 
			12'd1761 : q <= 23'h000000; 
			12'd1762 : q <= 23'h000000; 
			12'd1763 : q <= 23'h000000; 
			12'd1764 : q <= 23'h2530c2; 
			12'd1765 : q <= 23'h000000; 
			12'd1766 : q <= 23'h000000; 
			12'd1767 : q <= 23'h24bc43; 
			12'd1768 : q <= 23'h000000; 
			12'd1769 : q <= 23'h000000; 
			12'd1770 : q <= 23'h000000; 
			12'd1771 : q <= 23'h000000; 
			12'd1772 : q <= 23'h000000; 
			12'd1773 : q <= 23'h000000; 
			12'd1774 : q <= 23'h000000; 
			12'd1775 : q <= 23'h000000; 
			12'd1776 : q <= 23'h000000; 
			12'd1777 : q <= 23'h000000; 
			12'd1778 : q <= 23'h000000; 
			12'd1779 : q <= 23'h262021; 
			12'd1780 : q <= 23'h232021; 
			12'd1781 : q <= 23'h000000; 
			12'd1782 : q <= 23'h000000; 
			12'd1783 : q <= 23'h000000; 
			12'd1784 : q <= 23'h000000; 
			12'd1785 : q <= 23'h000000; 
			12'd1786 : q <= 23'h000000; 
			12'd1787 : q <= 23'h000000; 
			12'd1788 : q <= 23'h000000; 
			12'd1789 : q <= 23'h24a0a6; 
			12'd1790 : q <= 23'h000000; 
			12'd1791 : q <= 23'h000000; 
			12'd1792 : q <= 23'h000000; 
			12'd1793 : q <= 23'h000000; 
			12'd1794 : q <= 23'h241c41; 
			12'd1795 : q <= 23'h000000; 
			12'd1796 : q <= 23'h000000; 
			12'd1797 : q <= 23'h000000; 
			12'd1798 : q <= 23'h000000; 
			12'd1799 : q <= 23'h000000; 
			12'd1800 : q <= 23'h000000; 
			12'd1801 : q <= 23'h000000; 
			12'd1802 : q <= 23'h23c8a2; 
			12'd1803 : q <= 23'h22a4a3; 
			12'd1804 : q <= 23'h000000; 
			12'd1805 : q <= 23'h000000; 
			12'd1806 : q <= 23'h000000; 
			12'd1807 : q <= 23'h000000; 
			12'd1808 : q <= 23'h000000; 
			12'd1809 : q <= 23'h000000; 
			12'd1810 : q <= 23'h000000; 
			12'd1811 : q <= 23'h000000; 
			12'd1812 : q <= 23'h000000; 
			12'd1813 : q <= 23'h000000; 
			12'd1814 : q <= 23'h000000; 
			12'd1815 : q <= 23'h240c81; 
			12'd1816 : q <= 23'h000000; 
			12'd1817 : q <= 23'h000000; 
			12'd1818 : q <= 23'h000000; 
			12'd1819 : q <= 23'h000000; 
			12'd1820 : q <= 23'h000000; 
			12'd1821 : q <= 23'h274024; 
			12'd1822 : q <= 23'h000000; 
			12'd1823 : q <= 23'h274024; 
			12'd1824 : q <= 23'h251886; 
			12'd1825 : q <= 23'h000000; 
			12'd1826 : q <= 23'h000000; 
			12'd1827 : q <= 23'h26c463; 
			12'd1828 : q <= 23'h254941; 
			12'd1829 : q <= 23'h251823; 
			12'd1830 : q <= 23'h000000; 
			12'd1831 : q <= 23'h000000; 
			12'd1832 : q <= 23'h000000; 
			12'd1833 : q <= 23'h000000; 
			12'd1834 : q <= 23'h000000; 
			12'd1835 : q <= 23'h000000; 
			12'd1836 : q <= 23'h000000; 
			12'd1837 : q <= 23'h000000; 
			12'd1838 : q <= 23'h000000; 
			12'd1839 : q <= 23'h2444c3; 
			12'd1840 : q <= 23'h253d42; 
			12'd1841 : q <= 23'h2218e1; 
			12'd1842 : q <= 23'h2320a6; 
			12'd1843 : q <= 23'h000000; 
			12'd1844 : q <= 23'h000000; 
			12'd1845 : q <= 23'h000000; 
			12'd1846 : q <= 23'h23c041; 
			12'd1847 : q <= 23'h000000; 
			12'd1848 : q <= 23'h254842; 
			12'd1849 : q <= 23'h000000; 
			12'd1850 : q <= 23'h000000; 
			12'd1851 : q <= 23'h26c463; 
			12'd1852 : q <= 23'h000000; 
			12'd1853 : q <= 23'h26c463; 
			12'd1854 : q <= 23'h000000; 
			12'd1855 : q <= 23'h000000; 
			12'd1856 : q <= 23'h224463; 
			12'd1857 : q <= 23'h244443; 
			12'd1858 : q <= 23'h000000; 
			12'd1859 : q <= 23'h000000; 
			12'd1860 : q <= 23'h000000; 
			12'd1861 : q <= 23'h264443; 
			12'd1862 : q <= 23'h234443; 
			12'd1863 : q <= 23'h26c423; 
			12'd1864 : q <= 23'h234423; 
			12'd1865 : q <= 23'h000000; 
			12'd1866 : q <= 23'h000000; 
			12'd1867 : q <= 23'h000000; 
			12'd1868 : q <= 23'h000000; 
			12'd1869 : q <= 23'h000000; 
			12'd1870 : q <= 23'h000000; 
			12'd1871 : q <= 23'h26c064; 
			12'd1872 : q <= 23'h000000; 
			12'd1873 : q <= 23'h000000; 
			12'd1874 : q <= 23'h000000; 
			12'd1875 : q <= 23'h000000; 
			12'd1876 : q <= 23'h000000; 
			12'd1877 : q <= 23'h000000; 
			12'd1878 : q <= 23'h000000; 
			12'd1879 : q <= 23'h000000; 
			12'd1880 : q <= 23'h000000; 
			12'd1881 : q <= 23'h000000; 
			12'd1882 : q <= 23'h000000; 
			12'd1883 : q <= 23'h27c024; 
			12'd1884 : q <= 23'h000000; 
			12'd1885 : q <= 23'h24b861; 
			12'd1886 : q <= 23'h000000; 
			12'd1887 : q <= 23'h000000; 
			12'd1888 : q <= 23'h000000; 
			12'd1889 : q <= 23'h000000; 
			12'd1890 : q <= 23'h000000; 
			12'd1891 : q <= 23'h27c024; 
			12'd1892 : q <= 23'h224024; 
			12'd1893 : q <= 23'h000000; 
			12'd1894 : q <= 23'h000000; 
			12'd1895 : q <= 23'h2318a1; 
			12'd1896 : q <= 23'h000000; 
			12'd1897 : q <= 23'h000000; 
			12'd1898 : q <= 23'h22c421; 
			12'd1899 : q <= 23'h000000; 
			12'd1900 : q <= 23'h254941; 
			12'd1901 : q <= 23'h000000; 
			12'd1902 : q <= 23'h000000; 
			12'd1903 : q <= 23'h000000; 
			12'd1904 : q <= 23'h224c21; 
			12'd1905 : q <= 23'h000000; 
			12'd1906 : q <= 23'h000000; 
			12'd1907 : q <= 23'h000000; 
			12'd1908 : q <= 23'h253c61; 
			12'd1909 : q <= 23'h000000; 
			12'd1910 : q <= 23'h000000; 
			12'd1911 : q <= 23'h000000; 
			12'd1912 : q <= 23'h24c4e2; 
			12'd1913 : q <= 23'h21a0e1; 
			12'd1914 : q <= 23'h000000; 
			12'd1915 : q <= 23'h000000; 
			12'd1916 : q <= 23'h000000; 
			12'd1917 : q <= 23'h000000; 
			12'd1918 : q <= 23'h000000; 
			12'd1919 : q <= 23'h000000; 
			12'd1920 : q <= 23'h000000; 
			12'd1921 : q <= 23'h000000; 
			12'd1922 : q <= 23'h000000; 
			12'd1923 : q <= 23'h000000; 
			12'd1924 : q <= 23'h000000; 
			12'd1925 : q <= 23'h000000; 
			12'd1926 : q <= 23'h000000; 
			12'd1927 : q <= 23'h000000; 
			12'd1928 : q <= 23'h000000; 
			12'd1929 : q <= 23'h000000; 
			12'd1930 : q <= 23'h000000; 
			12'd1931 : q <= 23'h000000; 
			12'd1932 : q <= 23'h272c28; 
			12'd1933 : q <= 23'h000000; 
			12'd1934 : q <= 23'h000000; 
			12'd1935 : q <= 23'h244c41; 
			12'd1936 : q <= 23'h212505; 
			12'd1937 : q <= 23'h000000; 
			12'd1938 : q <= 23'h000000; 
			12'd1939 : q <= 23'h000000; 
			12'd1940 : q <= 23'h000000; 
			12'd1941 : q <= 23'h000000; 
			12'd1942 : q <= 23'h000000; 
			12'd1943 : q <= 23'h000000; 
			12'd1944 : q <= 23'h000000; 
			12'd1945 : q <= 23'h000000; 
			12'd1946 : q <= 23'h000000; 
			12'd1947 : q <= 23'h000000; 
			12'd1948 : q <= 23'h000000; 
			12'd1949 : q <= 23'h000000; 
			12'd1950 : q <= 23'h000000; 
			12'd1951 : q <= 23'h000000; 
			12'd1952 : q <= 23'h000000; 
			12'd1953 : q <= 23'h000000; 
			12'd1954 : q <= 23'h000000; 
			12'd1955 : q <= 23'h000000; 
			12'd1956 : q <= 23'h22a0a2; 
			12'd1957 : q <= 23'h000000; 
			12'd1958 : q <= 23'h253421; 
			12'd1959 : q <= 23'h000000; 
			12'd1960 : q <= 23'h000000; 
			12'd1961 : q <= 23'h000000; 
			12'd1962 : q <= 23'h000000; 
			12'd1963 : q <= 23'h000000; 
			12'd1964 : q <= 23'h000000; 
			12'd1965 : q <= 23'h000000; 
			12'd1966 : q <= 23'h000000; 
			12'd1967 : q <= 23'h000000; 
			12'd1968 : q <= 23'h000000; 
			12'd1969 : q <= 23'h000000; 
			12'd1970 : q <= 23'h233484; 
			12'd1971 : q <= 23'h24bc43; 
			12'd1972 : q <= 23'h000000; 
			12'd1973 : q <= 23'h253025; 
			12'd1974 : q <= 23'h000000; 
			12'd1975 : q <= 23'h000000; 
			12'd1976 : q <= 23'h000000; 
			12'd1977 : q <= 23'h224463; 
			12'd1978 : q <= 23'h000000; 
			12'd1979 : q <= 23'h000000; 
			12'd1980 : q <= 23'h000000; 
			12'd1981 : q <= 23'h000000; 
			12'd1982 : q <= 23'h000000; 
			12'd1983 : q <= 23'h000000; 
			12'd1984 : q <= 23'h000000; 
			12'd1985 : q <= 23'h000000; 
			12'd1986 : q <= 23'h000000; 
			12'd1987 : q <= 23'h000000; 
			12'd1988 : q <= 23'h25b421; 
			12'd1989 : q <= 23'h243421; 
			12'd1990 : q <= 23'h000000; 
			12'd1991 : q <= 23'h000000; 
			12'd1992 : q <= 23'h000000; 
			12'd1993 : q <= 23'h000000; 
			12'd1994 : q <= 23'h000000; 
			12'd1995 : q <= 23'h000000; 
			12'd1996 : q <= 23'h000000; 
			12'd1997 : q <= 23'h000000; 
			12'd1998 : q <= 23'h2240c2; 
			12'd1999 : q <= 23'h000000; 
			12'd2000 : q <= 23'h000000; 
			12'd2001 : q <= 23'h253844; 
			12'd2002 : q <= 23'h000000; 
			12'd2003 : q <= 23'h000000; 
			12'd2004 : q <= 23'h000000; 
			12'd2005 : q <= 23'h000000; 
			12'd2006 : q <= 23'h000000; 
			12'd2007 : q <= 23'h219825; 
			12'd2008 : q <= 23'h000000; 
			12'd2009 : q <= 23'h000000; 
			12'd2010 : q <= 23'h000000; 
			12'd2011 : q <= 23'h000000; 
			12'd2012 : q <= 23'h269861; 
			12'd2013 : q <= 23'h000000; 
			12'd2014 : q <= 23'h000000; 
			12'd2015 : q <= 23'h000000; 
			12'd2016 : q <= 23'h000000; 
			12'd2017 : q <= 23'h000000; 
			12'd2018 : q <= 23'h000000; 
			12'd2019 : q <= 23'h000000; 
			12'd2020 : q <= 23'h000000; 
			12'd2021 : q <= 23'h000000; 
			12'd2022 : q <= 23'h000000; 
			12'd2023 : q <= 23'h000000; 
			12'd2024 : q <= 23'h000000; 
			12'd2025 : q <= 23'h253903; 
			12'd2026 : q <= 23'h262021; 
			12'd2027 : q <= 23'h000000; 
			12'd2028 : q <= 23'h000000; 
			12'd2029 : q <= 23'h000000; 
			12'd2030 : q <= 23'h000000; 
			12'd2031 : q <= 23'h000000; 
			12'd2032 : q <= 23'h000000; 
			12'd2033 : q <= 23'h000000; 
			12'd2034 : q <= 23'h000000; 
			12'd2035 : q <= 23'h000000; 
			12'd2036 : q <= 23'h24c423; 
			12'd2037 : q <= 23'h000000; 
			12'd2038 : q <= 23'h000000; 
			12'd2039 : q <= 23'h000000; 
			12'd2040 : q <= 23'h000000; 
			12'd2041 : q <= 23'h000000; 
			12'd2042 : q <= 23'h000000; 
			12'd2043 : q <= 23'h232021; 
			12'd2044 : q <= 23'h000000; 
			12'd2045 : q <= 23'h000000; 
			12'd2046 : q <= 23'h000000; 
			12'd2047 : q <= 23'h20ac28; 
			12'd2048 : q <= 23'h000000; 
			12'd2049 : q <= 23'h000000; 
			12'd2050 : q <= 23'h000000; 
			12'd2051 : q <= 23'h000000; 
			12'd2052 : q <= 23'h000000; 
			12'd2053 : q <= 23'h000000; 
			12'd2054 : q <= 23'h000000; 
			12'd2055 : q <= 23'h000000; 
			12'd2056 : q <= 23'h000000; 
			12'd2057 : q <= 23'h249123; 
			12'd2058 : q <= 23'h000000; 
			12'd2059 : q <= 23'h000000; 
			12'd2060 : q <= 23'h000000; 
			12'd2061 : q <= 23'h000000; 
			12'd2062 : q <= 23'h000000; 
			12'd2063 : q <= 23'h000000; 
			12'd2064 : q <= 23'h000000; 
			12'd2065 : q <= 23'h000000; 
			12'd2066 : q <= 23'h000000; 
			12'd2067 : q <= 23'h000000; 
			12'd2068 : q <= 23'h000000; 
			12'd2069 : q <= 23'h000000; 
			12'd2070 : q <= 23'h268862; 
			12'd2071 : q <= 23'h000000; 
			12'd2072 : q <= 23'h000000; 
			12'd2073 : q <= 23'h000000; 
			12'd2074 : q <= 23'h000000; 
			12'd2075 : q <= 23'h000000; 
			12'd2076 : q <= 23'h000000; 
			12'd2077 : q <= 23'h000000; 
			12'd2078 : q <= 23'h000000; 
			12'd2079 : q <= 23'h000000; 
			12'd2080 : q <= 23'h000000; 
			12'd2081 : q <= 23'h000000; 
			12'd2082 : q <= 23'h000000; 
			12'd2083 : q <= 23'h241841; 
			12'd2084 : q <= 23'h000000; 
			12'd2085 : q <= 23'h000000; 
			12'd2086 : q <= 23'h000000; 
			12'd2087 : q <= 23'h000000; 
			12'd2088 : q <= 23'h000000; 
			12'd2089 : q <= 23'h220862; 
			12'd2090 : q <= 23'h000000; 
			12'd2091 : q <= 23'h000000; 
			12'd2092 : q <= 23'h000000; 
			12'd2093 : q <= 23'h000000; 
			12'd2094 : q <= 23'h000000; 
			12'd2095 : q <= 23'h000000; 
			12'd2096 : q <= 23'h243046; 
			12'd2097 : q <= 23'h000000; 
			12'd2098 : q <= 23'h000000; 
			12'd2099 : q <= 23'h000000; 
			12'd2100 : q <= 23'h000000; 
			12'd2101 : q <= 23'h000000; 
			12'd2102 : q <= 23'h000000; 
			12'd2103 : q <= 23'h24c042; 
			12'd2104 : q <= 23'h26c443; 
			12'd2105 : q <= 23'h000000; 
			12'd2106 : q <= 23'h281024; 
			12'd2107 : q <= 23'h219024; 
			12'd2108 : q <= 23'h000000; 
			12'd2109 : q <= 23'h000000; 
			12'd2110 : q <= 23'h000000; 
			12'd2111 : q <= 23'h000000; 
			12'd2112 : q <= 23'h000000; 
			12'd2113 : q <= 23'h000000; 
			12'd2114 : q <= 23'h000000; 
			12'd2115 : q <= 23'h000000; 
			12'd2116 : q <= 23'h000000; 
			12'd2117 : q <= 23'h000000; 
			12'd2118 : q <= 23'h000000; 
			12'd2119 : q <= 23'h000000; 
			12'd2120 : q <= 23'h000000; 
			12'd2121 : q <= 23'h000000; 
			12'd2122 : q <= 23'h000000; 
			12'd2123 : q <= 23'h000000; 
			12'd2124 : q <= 23'h000000; 
			12'd2125 : q <= 23'h000000; 
			12'd2126 : q <= 23'h000000; 
			12'd2127 : q <= 23'h000000; 
			12'd2128 : q <= 23'h000000; 
			12'd2129 : q <= 23'h000000; 
			12'd2130 : q <= 23'h000000; 
			12'd2131 : q <= 23'h000000; 
			12'd2132 : q <= 23'h000000; 
			12'd2133 : q <= 23'h000000; 
			12'd2134 : q <= 23'h000000; 
			12'd2135 : q <= 23'h228ca3;
			default	 : q <= 23'h000000;
		endcase	
	end
	assign out = q;
endmodule