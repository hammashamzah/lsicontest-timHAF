module nnodes_stagethreshold_rom(
	input clk,
	input [4:0] addr,
	output[23:0] out
);
	reg[23:0] q;

	always @(posedge clk)
	begin
		case(addr)
			12'd1   : q <= 24'd196818;
			12'd2   : q <= 24'd1050356;
			12'd3   : q <= 24'd1378687;
			12'd4   : q <= 24'd2560617;
			12'd5   : q <= 24'd2166610;
			12'd6   : q <= 24'd2888962;
			12'd7   : q <= 24'd3282923;
			12'd8   : q <= 24'd3348615;
			12'd9   : q <= 24'd3676967;
			12'd10	: q <= 24'd4661901;
			12'd11	: q <= 24'd5252891;
			12'd12	: q <= 24'd6763164;
			12'd13	: q <= 24'd7288478;
			12'd14	: q <= 24'd6697515;
			12'd15	: q <= 24'd8864427;
			12'd16	: q <= 24'd8995762;
			12'd17	: q <= 24'd9192762;
			12'd18	: q <= 24'd10506047;
			12'd19	: q <= 24'd11622322;
			12'd20	: q <= 24'd11950656;
			12'd21	: q <= 24'd13854911;
			12'd22	: q <= 24'd13986242;
			default	: q <= 24'd00000000;
		endcase	
	end
	assign out = q;
endmodule