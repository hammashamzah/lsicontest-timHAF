module nnodes_left_right_rom(
	input clk,
	input [11:0] addr,
	output[27:0] out
);
	reg[27:0] q;

	always @(posedge clk)
	begin
		case(addr)
			12'd1    : q <= 28'h00108d6;
			12'd2    : q <= 28'h00326bf;
			12'd3    : q <= 28'h00117a3;
			12'd4    : q <= 28'h00011b6;
			12'd5    : q <= 28'h0002daa;
			12'd6    : q <= 28'h0012ba7;
			12'd7    : q <= 28'h0029617;
			12'd8    : q <= 28'h000249a;
			12'd9    : q <= 28'h0095eca;
			12'd10   : q <= 28'h0029d35;
			12'd11   : q <= 28'h00248a2;
			12'd12   : q <= 28'h0003894;
			12'd13   : q <= 28'h0003d94;
			12'd14   : q <= 28'h0008e22;
			12'd15   : q <= 28'hfe8d978;
			12'd16   : q <= 28'h0009948;
			12'd17   : q <= 28'h0126fb4;
			12'd18   : q <= 28'h0004d9a;
			12'd19   : q <= 28'hfff2e91;
			12'd20   : q <= 28'hffcaa24;
			12'd21   : q <= 28'h000a120;
			12'd22   : q <= 28'h0001f9e;
			12'd23   : q <= 28'h0002491;
			12'd24   : q <= 28'h0002a97;
			12'd25   : q <= 28'h0004592;
			12'd26   : q <= 28'hfff3094;
			12'd27   : q <= 28'h0003b91;
			12'd28   : q <= 28'h0004698;
			12'd29   : q <= 28'hffe2c8d;
			12'd30   : q <= 28'hffd228e;
			12'd31   : q <= 28'h0015c9e;
			12'd32   : q <= 28'hfec178c;
			12'd33   : q <= 28'h0005f92;
			12'd34   : q <= 28'h0009854;
			12'd35   : q <= 28'hff32f8f;
			12'd36   : q <= 28'h0005c9c;
			12'd37   : q <= 28'h0009958;
			12'd38   : q <= 28'h0016ab2;
			12'd39   : q <= 28'h00173c7;
			12'd40   : q <= 28'h0068b21;
			12'd41   : q <= 28'h000249e;
			12'd42   : q <= 28'h0009e30;
			12'd43   : q <= 28'h0002695;
			12'd44   : q <= 28'h00146a2;
			12'd45   : q <= 28'h0019637;
			12'd46   : q <= 28'h000964c;
			12'd47   : q <= 28'h0003c96;
			12'd48   : q <= 28'hffb1f84;
			12'd49   : q <= 28'hfff4394;
			12'd50   : q <= 28'h0005d91;
			12'd51   : q <= 28'h00d6ec1;
			12'd52   : q <= 28'h000368f;
			12'd53   : q <= 28'h0009043;
			12'd54   : q <= 28'h0069446;
			12'd55   : q <= 28'h0004593;
			12'd56   : q <= 28'h0008b3b;
			12'd57   : q <= 28'h0008834;
			12'd58   : q <= 28'h0008a4e;
			12'd59   : q <= 28'h0005e9c;
			12'd60   : q <= 28'h0005b9a;
			12'd61   : q <= 28'h0003089;
			12'd62   : q <= 28'h000628d;
			12'd63   : q <= 28'h0006eb5;
			12'd64   : q <= 28'h00066a3;
			12'd65   : q <= 28'hffd3c8b;
			12'd66   : q <= 28'h0019452;
			12'd67   : q <= 28'h0008d4a;
			12'd68   : q <= 28'hfff2d85;
			12'd69   : q <= 28'h0004d8d;
			12'd70   : q <= 28'h00571b2;
			12'd71   : q <= 28'h000478c;
			12'd72   : q <= 28'h001863d;
			12'd73   : q <= 28'h0006eb2;
			12'd74   : q <= 28'hfff4e8a;
			12'd75   : q <= 28'h0008d4f;
			12'd76   : q <= 28'h0078a2d;
			12'd77   : q <= 28'h002841f;
			12'd78   : q <= 28'h0058754;
			12'd79   : q <= 28'hffebf71;
			12'd80   : q <= 28'h000349b;
			12'd81   : q <= 28'h0009520;
			12'd82   : q <= 28'h0001892;
			12'd83   : q <= 28'h0002d91;
			12'd84   : q <= 28'h0002994;
			12'd85   : q <= 28'h000358d;
			12'd86   : q <= 28'h000912f;
			12'd87   : q <= 28'h0028238;
			12'd88   : q <= 28'hff0b667;
			12'd89   : q <= 28'hffe418b;
			12'd90   : q <= 28'h0002b8f;
			12'd91   : q <= 28'h0008a43;
			12'd92   : q <= 28'h0045fa7;
			12'd93   : q <= 28'hfff438d;
			12'd94   : q <= 28'hffd338d;
			12'd95   : q <= 28'h0008f4d;
			12'd96   : q <= 28'h0004590;
			12'd97   : q <= 28'hfff238b;
			12'd98   : q <= 28'h0002d8b;
			12'd99   : q <= 28'hffe9247;
			12'd100  : q <= 28'hfff3c8c; 
			12'd101  : q <= 28'h0018f54; 
			12'd102  : q <= 28'hfff2989; 
			12'd103  : q <= 28'h003853a; 
			12'd104  : q <= 28'hffeb36c; 
			12'd105  : q <= 28'hffe4689; 
			12'd106  : q <= 28'h0296fbe; 
			12'd107  : q <= 28'h0019242; 
			12'd108  : q <= 28'h0003589; 
			12'd109  : q <= 28'hffdc274; 
			12'd110  : q <= 28'hff02088; 
			12'd111  : q <= 28'h002548f; 
			12'd112  : q <= 28'h0058c46; 
			12'd113  : q <= 28'h0002d9d; 
			12'd114  : q <= 28'h0009c2e; 
			12'd115  : q <= 28'h0001992; 
			12'd116  : q <= 28'h0008e3c; 
			12'd117  : q <= 28'h0003995; 
			12'd118  : q <= 28'h0004394; 
			12'd119  : q <= 28'h001943f; 
			12'd120  : q <= 28'hffd2e8c; 
			12'd121  : q <= 28'h000569a; 
			12'd122  : q <= 28'h0003a8b; 
			12'd123  : q <= 28'h000903d; 
			12'd124  : q <= 28'h0006498; 
			12'd125  : q <= 28'h0078628; 
			12'd126  : q <= 28'h0096bac; 
			12'd127  : q <= 28'hffa308c; 
			12'd128  : q <= 28'hfff2285; 
			12'd129  : q <= 28'h000609c; 
			12'd130  : q <= 28'hffb448a; 
			12'd131  : q <= 28'h0018939; 
			12'd132  : q <= 28'h011893e; 
			12'd133  : q <= 28'h0003d89; 
			12'd134  : q <= 28'h0008a50; 
			12'd135  : q <= 28'h0056aa8; 
			12'd136  : q <= 28'h000478c; 
			12'd137  : q <= 28'h0008630; 
			12'd138  : q <= 28'h0009155; 
			12'd139  : q <= 28'h003883d; 
			12'd140  : q <= 28'hfff9966; 
			12'd141  : q <= 28'hff2d174; 
			12'd142  : q <= 28'hfff3889; 
			12'd143  : q <= 28'h00170b7; 
			12'd144  : q <= 28'h0018c47; 
			12'd145  : q <= 28'h000a266; 
			12'd146  : q <= 28'h0005987; 
			12'd147  : q <= 28'hfff1c85; 
			12'd148  : q <= 28'hff33d8b; 
			12'd149  : q <= 28'hffec271; 
			12'd150  : q <= 28'h000418c; 
			12'd151  : q <= 28'h000ac6c; 
			12'd152  : q <= 28'h0048c3a; 
			12'd153  : q <= 28'h0009c66; 
			12'd154  : q <= 28'h0018727; 
			12'd155  : q <= 28'hfff2c86; 
			12'd156  : q <= 28'hffda86e; 
			12'd157  : q <= 28'hfff9c25; 
			12'd158  : q <= 28'h0004396; 
			12'd159  : q <= 28'h004962d; 
			12'd160  : q <= 28'h000288f; 
			12'd161  : q <= 28'h0003092; 
			12'd162  : q <= 28'h0004a8f; 
			12'd163  : q <= 28'hfe73190; 
			12'd164  : q <= 28'h000508c; 
			12'd165  : q <= 28'hffd4093; 
			12'd166  : q <= 28'h001935d; 
			12'd167  : q <= 28'h0004897; 
			12'd168  : q <= 28'h001679e; 
			12'd169  : q <= 28'h0009450; 
			12'd170  : q <= 28'h00d8d31; 
			12'd171  : q <= 28'h00367aa; 
			12'd172  : q <= 28'h0005a92; 
			12'd173  : q <= 28'h0004d8f; 
			12'd174  : q <= 28'hfffb775; 
			12'd175  : q <= 28'h0008f4b; 
			12'd176  : q <= 28'h00176c3; 
			12'd177  : q <= 28'h003882d; 
			12'd178  : q <= 28'hff22b88; 
			12'd179  : q <= 28'h000619a; 
			12'd180  : q <= 28'hffe2688; 
			12'd181  : q <= 28'hffe3588; 
			12'd182  : q <= 28'h0006885; 
			12'd183  : q <= 28'h0009159; 
			12'd184  : q <= 28'h0038839; 
			12'd185  : q <= 28'hffa2785; 
			12'd186  : q <= 28'h0008c61; 
			12'd187  : q <= 28'h0006ca9; 
			12'd188  : q <= 28'hffb3789; 
			12'd189  : q <= 28'h000aa6b; 
			12'd190  : q <= 28'hfff3a89; 
			12'd191  : q <= 28'h0006eaf; 
			12'd192  : q <= 28'h0039558; 
			12'd193  : q <= 28'h000b36e; 
			12'd194  : q <= 28'h0004a85; 
			12'd195  : q <= 28'h0004c8c; 
			12'd196  : q <= 28'h0027dd1; 
			12'd197  : q <= 28'hffc2586; 
			12'd198  : q <= 28'h0047abc; 
			12'd199  : q <= 28'h000bc72; 
			12'd200  : q <= 28'hffe598d; 
			12'd201  : q <= 28'hffd3c88; 
			12'd202  : q <= 28'hffa3283; 
			12'd203  : q <= 28'h0008f56; 
			12'd204  : q <= 28'hfea1084; 
			12'd205  : q <= 28'h000bb72; 
			12'd206  : q <= 28'h0006999; 
			12'd207  : q <= 28'h00044aa; 
			12'd208  : q <= 28'h0009d40; 
			12'd209  : q <= 28'h000933d; 
			12'd210  : q <= 28'h0009140; 
			12'd211  : q <= 28'hfff2a8e; 
			12'd212  : q <= 28'hff59c79; 
			12'd213  : q <= 28'h0009248; 
			12'd214  : q <= 28'h0036899; 
			12'd215  : q <= 28'h0009245; 
			12'd216  : q <= 28'h0018653; 
			12'd217  : q <= 28'h000af6b; 
			12'd218  : q <= 28'hfff538b; 
			12'd219  : q <= 28'h0018b3b; 
			12'd220  : q <= 28'h0008e45; 
			12'd221  : q <= 28'h0005e96; 
			12'd222  : q <= 28'hfed368a; 
			12'd223  : q <= 28'h0048d45; 
			12'd224  : q <= 28'h000659a; 
			12'd225  : q <= 28'h0078624; 
			12'd226  : q <= 28'h0005697; 
			12'd227  : q <= 28'h0008c4d; 
			12'd228  : q <= 28'h000568d; 
			12'd229  : q <= 28'h0009056; 
			12'd230  : q <= 28'hfe61085; 
			12'd231  : q <= 28'h009831a; 
			12'd232  : q <= 28'h000638e; 
			12'd233  : q <= 28'h0058630; 
			12'd234  : q <= 28'h000aa77; 
			12'd235  : q <= 28'h000b76e; 
			12'd236  : q <= 28'h0004d90; 
			12'd237  : q <= 28'hfff2e86; 
			12'd238  : q <= 28'h000568b; 
			12'd239  : q <= 28'h00068a0; 
			12'd240  : q <= 28'hffe5691; 
			12'd241  : q <= 28'h0006ba6; 
			12'd242  : q <= 28'hfff428a; 
			12'd243  : q <= 28'h0009d65; 
			12'd244  : q <= 28'hffe2985; 
			12'd245  : q <= 28'h000518c; 
			12'd246  : q <= 28'h003699c; 
			12'd247  : q <= 28'hffb1a85; 
			12'd248  : q <= 28'hfe0d97d; 
			12'd249  : q <= 28'h000508c; 
			12'd250  : q <= 28'h0147c9b; 
			12'd251  : q <= 28'hfecd676; 
			12'd252  : q <= 28'hfff3087; 
			12'd253  : q <= 28'h0008642; 
			12'd254  : q <= 28'h0006c92; 
			12'd255  : q <= 28'h000b173; 
			12'd256  : q <= 28'h0029769; 
			12'd257  : q <= 28'h000a56e; 
			12'd258  : q <= 28'hffe9d3f; 
			12'd259  : q <= 28'h000923b; 
			12'd260  : q <= 28'h0003694; 
			12'd261  : q <= 28'h0014b96; 
			12'd262  : q <= 28'h0004c94; 
			12'd263  : q <= 28'hffe4890; 
			12'd264  : q <= 28'h0025a9b; 
			12'd265  : q <= 28'h0008f45; 
			12'd266  : q <= 28'h000995d; 
			12'd267  : q <= 28'h000468b; 
			12'd268  : q <= 28'h0016eb4; 
			12'd269  : q <= 28'hff23f87; 
			12'd270  : q <= 28'h0018c3f; 
			12'd271  : q <= 28'h0006492; 
			12'd272  : q <= 28'h00170bd; 
			12'd273  : q <= 28'h0018b3f; 
			12'd274  : q <= 28'h0004188; 
			12'd275  : q <= 28'hfff4588; 
			12'd276  : q <= 28'h000518d; 
			12'd277  : q <= 28'h0006da7; 
			12'd278  : q <= 28'h0009761; 
			12'd279  : q <= 28'h0016192; 
			12'd280  : q <= 28'h0002c86; 
			12'd281  : q <= 28'h0005c92; 
			12'd282  : q <= 28'h0008a4d; 
			12'd283  : q <= 28'hffd528e; 
			12'd284  : q <= 28'h0066ea6; 
			12'd285  : q <= 28'h0005b8f; 
			12'd286  : q <= 28'h000598e; 
			12'd287  : q <= 28'hffd2d88; 
			12'd288  : q <= 28'h0009d6c; 
			12'd289  : q <= 28'h0048a37; 
			12'd290  : q <= 28'h000a56f; 
			12'd291  : q <= 28'h0008a5a; 
			12'd292  : q <= 28'hfff4788; 
			12'd293  : q <= 28'h001915e; 
			12'd294  : q <= 28'hffec675; 
			12'd295  : q <= 28'h0008866; 
			12'd296  : q <= 28'h0008f60; 
			12'd297  : q <= 28'hffe4a84; 
			12'd298  : q <= 28'h0008d5e; 
			12'd299  : q <= 28'hfff6091; 
			12'd300  : q <= 28'hfffb372; 
			12'd301  : q <= 28'hfff3b88; 
			12'd302  : q <= 28'h0009669; 
			12'd303  : q <= 28'h0005f8f; 
			12'd304  : q <= 28'h00a8745; 
			12'd305  : q <= 28'h00178ab; 
			12'd306  : q <= 28'h0018429; 
			12'd307  : q <= 28'h0018a4b; 
			12'd308  : q <= 28'hffdb574; 
			12'd309  : q <= 28'h007855b; 
			12'd310  : q <= 28'h000598b; 
			12'd311  : q <= 28'h0009667; 
			12'd312  : q <= 28'hffeac71; 
			12'd313  : q <= 28'h004872e; 
			12'd314  : q <= 28'hfff9743; 
			12'd315  : q <= 28'h0003b92; 
			12'd316  : q <= 28'hffe2a90; 
			12'd317  : q <= 28'h0158a32; 
			12'd318  : q <= 28'h0005799; 
			12'd319  : q <= 28'h0015f9b; 
			12'd320  : q <= 28'h000418e; 
			12'd321  : q <= 28'h0004b8d; 
			12'd322  : q <= 28'hffec172; 
			12'd323  : q <= 28'h0088e44; 
			12'd324  : q <= 28'h000904c; 
			12'd325  : q <= 28'hffa4682; 
			12'd326  : q <= 28'h0008e4f; 
			12'd327  : q <= 28'h0005591; 
			12'd328  : q <= 28'h0004c88; 
			12'd329  : q <= 28'hfde258a; 
			12'd330  : q <= 28'h0005f91; 
			12'd331  : q <= 28'hff6468c; 
			12'd332  : q <= 28'h0005f93; 
			12'd333  : q <= 28'hfffc079; 
			12'd334  : q <= 28'h0008a4b; 
			12'd335  : q <= 28'h0009d6d; 
			12'd336  : q <= 28'h0003485; 
			12'd337  : q <= 28'h007862a; 
			12'd338  : q <= 28'h0008647; 
			12'd339  : q <= 28'hffeb27b; 
			12'd340  : q <= 28'h0016da2; 
			12'd341  : q <= 28'h0004b89; 
			12'd342  : q <= 28'h00173bd; 
			12'd343  : q <= 28'hffe508a; 
			12'd344  : q <= 28'h0068321; 
			12'd345  : q <= 28'h0098442; 
			12'd346  : q <= 28'h0058328; 
			12'd347  : q <= 28'h0008e70; 
			12'd348  : q <= 28'h0008e5e; 
			12'd349  : q <= 28'h000568e; 
			12'd350  : q <= 28'h0008957; 
			12'd351  : q <= 28'hfff9c6f; 
			12'd352  : q <= 28'hff43c84; 
			12'd353  : q <= 28'hff7bb79; 
			12'd354  : q <= 28'h0008a57; 
			12'd355  : q <= 28'h000488e; 
			12'd356  : q <= 28'hfece978; 
			12'd357  : q <= 28'h0009a65; 
			12'd358  : q <= 28'h0008f62; 
			12'd359  : q <= 28'hfef3987; 
			12'd360  : q <= 28'h0036895; 
			12'd361  : q <= 28'hfff4886; 
			12'd362  : q <= 28'h009811a; 
			12'd363  : q <= 28'h0009d6f; 
			12'd364  : q <= 28'h00273c2; 
			12'd365  : q <= 28'h001862f; 
			12'd366  : q <= 28'h004853b; 
			12'd367  : q <= 28'h0048b53; 
			12'd368  : q <= 28'hff7b374; 
			12'd369  : q <= 28'hffb438a; 
			12'd370  : q <= 28'h00172b6; 
			12'd371  : q <= 28'h0006c8c; 
			12'd372  : q <= 28'h0008850; 
			12'd373  : q <= 28'h0088357; 
			12'd374  : q <= 28'h0005a8b; 
			12'd375  : q <= 28'hffe4888; 
			12'd376  : q <= 28'hfffb073; 
			12'd377  : q <= 28'hffe2b85; 
			12'd378  : q <= 28'h000874c; 
			12'd379  : q <= 28'h000a672; 
			12'd380  : q <= 28'h0005389; 
			12'd381  : q <= 28'hffac07a; 
			12'd382  : q <= 28'h0018853; 
			12'd383  : q <= 28'h0027592; 
			12'd384  : q <= 28'hffe4285; 
			12'd385  : q <= 28'h00153af; 
			12'd386  : q <= 28'h0009540; 
			12'd387  : q <= 28'h0009247; 
			12'd388  : q <= 28'h002408d; 
			12'd389  : q <= 28'h0003d8b; 
			12'd390  : q <= 28'h002659f; 
			12'd391  : q <= 28'h000904c; 
			12'd392  : q <= 28'hfff378a; 
			12'd393  : q <= 28'h0003c89; 
			12'd394  : q <= 28'h0006192; 
			12'd395  : q <= 28'h0004086; 
			12'd396  : q <= 28'h0009962; 
			12'd397  : q <= 28'h000915d; 
			12'd398  : q <= 28'hff92689; 
			12'd399  : q <= 28'h0005e8e; 
			12'd400  : q <= 28'hfffad74; 
			12'd401  : q <= 28'h000894b; 
			12'd402  : q <= 28'hffc2a88; 
			12'd403  : q <= 28'hfff3283; 
			12'd404  : q <= 28'h00177b3; 
			12'd405  : q <= 28'hff81d82; 
			12'd406  : q <= 28'h0178321; 
			12'd407  : q <= 28'h0005c8b; 
			12'd408  : q <= 28'h0037dc4; 
			12'd409  : q <= 28'h0008952; 
			12'd410  : q <= 28'hff42f85; 
			12'd411  : q <= 28'h000628d; 
			12'd412  : q <= 28'h0026d9c; 
			12'd413  : q <= 28'h0004a87; 
			12'd414  : q <= 28'hff6c17c; 
			12'd415  : q <= 28'hffa4886; 
			12'd416  : q <= 28'h00a7ca0; 
			12'd417  : q <= 28'hffab575; 
			12'd418  : q <= 28'h000678c; 
			12'd419  : q <= 28'h00573ad; 
			12'd420  : q <= 28'h0038b61; 
			12'd421  : q <= 28'h0006b96; 
			12'd422  : q <= 28'hffe618e; 
			12'd423  : q <= 28'hfffb975; 
			12'd424  : q <= 28'h0007897; 
			12'd425  : q <= 28'h022832e; 
			12'd426  : q <= 28'h0008a5f; 
			12'd427  : q <= 28'h0003d83; 
			12'd428  : q <= 28'hfffa879; 
			12'd429  : q <= 28'h0006ba1; 
			12'd430  : q <= 28'h0008d5e; 
			12'd431  : q <= 28'hffa2b82; 
			12'd432  : q <= 28'hff93084; 
			12'd433  : q <= 28'h00071a1; 
			12'd434  : q <= 28'hff73f89; 
			12'd435  : q <= 28'h000895d; 
			12'd436  : q <= 28'h0008d5a; 
			12'd437  : q <= 28'h0006991; 
			12'd438  : q <= 28'hfff1985; 
			12'd439  : q <= 28'hffa1780; 
			12'd440  : q <= 28'h001799f; 
			12'd441  : q <= 28'hfff3783; 
			12'd442  : q <= 28'h0008a5f; 
			12'd443  : q <= 28'hffcc777; 
			12'd444  : q <= 28'h0008c6c; 
			12'd445  : q <= 28'h0008859; 
			12'd446  : q <= 28'hffeb179; 
			12'd447  : q <= 28'h00c8113; 
			12'd448  : q <= 28'h000608d; 
			12'd449  : q <= 28'h0004e89; 
			12'd450  : q <= 28'h000a977; 
			12'd451  : q <= 28'h000a86f; 
			12'd452  : q <= 28'h002853b; 
			12'd453  : q <= 28'h000854c; 
			12'd454  : q <= 28'hff7b97c; 
			12'd455  : q <= 28'h0004f85; 
			12'd456  : q <= 28'h0005085; 
			12'd457  : q <= 28'h00074a8; 
			12'd458  : q <= 28'hff42e85; 
			12'd459  : q <= 28'h000b977; 
			12'd460  : q <= 28'h0007097; 
			12'd461  : q <= 28'h0005989; 
			12'd462  : q <= 28'h0047dd4; 
			12'd463  : q <= 28'h0005b89; 
			12'd464  : q <= 28'h0006f98; 
			12'd465  : q <= 28'hffe9d4e; 
			12'd466  : q <= 28'h0009450; 
			12'd467  : q <= 28'h0004191; 
			12'd468  : q <= 28'h0005e97; 
			12'd469  : q <= 28'h0003b8c; 
			12'd470  : q <= 28'h0005391; 
			12'd471  : q <= 28'h0005f95; 
			12'd472  : q <= 28'h000578d; 
			12'd473  : q <= 28'h0004789; 
			12'd474  : q <= 28'h000428c; 
			12'd475  : q <= 28'h0006aa1; 
			12'd476  : q <= 28'h0009667; 
			12'd477  : q <= 28'h002853b; 
			12'd478  : q <= 28'hffc4686; 
			12'd479  : q <= 28'h000925e; 
			12'd480  : q <= 28'h000728d; 
			12'd481  : q <= 28'h0004887; 
			12'd482  : q <= 28'h0017094; 
			12'd483  : q <= 28'hffd4c87; 
			12'd484  : q <= 28'hffdc579; 
			12'd485  : q <= 28'h0005f8e; 
			12'd486  : q <= 28'hffe5c87; 
			12'd487  : q <= 28'h0008959; 
			12'd488  : q <= 28'hfffb177; 
			12'd489  : q <= 28'hffdc577; 
			12'd490  : q <= 28'hffe5688; 
			12'd491  : q <= 28'h0008854; 
			12'd492  : q <= 28'hffdaf79; 
			12'd493  : q <= 28'h0005b89; 
			12'd494  : q <= 28'h0008d5a; 
			12'd495  : q <= 28'h0018120; 
			12'd496  : q <= 28'h0078629; 
			12'd497  : q <= 28'hfffb675; 
			12'd498  : q <= 28'h0008a59; 
			12'd499  : q <= 28'hfeb3e84; 
			12'd500  : q <= 28'h0006393; 
			12'd501  : q <= 28'h0005688; 
			12'd502  : q <= 28'h00075a3; 
			12'd503  : q <= 28'h0009369; 
			12'd504  : q <= 28'h0037cb5; 
			12'd505  : q <= 28'h000864a; 
			12'd506  : q <= 28'hff92685; 
			12'd507  : q <= 28'hff9067f; 
			12'd508  : q <= 28'h0008b67; 
			12'd509  : q <= 28'h0016d96; 
			12'd510  : q <= 28'hfeeaf7d; 
			12'd511  : q <= 28'hffc5688; 
			12'd512  : q <= 28'h003769c; 
			12'd513  : q <= 28'h0028857; 
			12'd514  : q <= 28'h0007695; 
			12'd515  : q <= 28'h0008549; 
			12'd516  : q <= 28'h0007b98; 
			12'd517  : q <= 28'hfffe479; 
			12'd518  : q <= 28'hfff3488; 
			12'd519  : q <= 28'h00075ac; 
			12'd520  : q <= 28'h0018648; 
			12'd521  : q <= 28'h0006992; 
			12'd522  : q <= 28'h0028547; 
			12'd523  : q <= 28'h0008654; 
			12'd524  : q <= 28'h00073a0; 
			12'd525  : q <= 28'h0068333; 
			12'd526  : q <= 28'hffec77c; 
			12'd527  : q <= 28'h0006d96; 
			12'd528  : q <= 28'hfff5a87; 
			12'd529  : q <= 28'hfffaf75; 
			12'd530  : q <= 28'h0005b8c; 
			12'd531  : q <= 28'h0005686; 
			12'd532  : q <= 28'h000578b; 
			12'd533  : q <= 28'hffea772; 
			12'd534  : q <= 28'h0008764; 
			12'd535  : q <= 28'hff9af75; 
			12'd536  : q <= 28'h0006789; 
			12'd537  : q <= 28'h0008a5e; 
			12'd538  : q <= 28'h00077a5; 
			12'd539  : q <= 28'h0009768; 
			12'd540  : q <= 28'hffd5d87; 
			12'd541  : q <= 28'hffc4483; 
			12'd542  : q <= 28'hfffad7c; 
			12'd543  : q <= 28'h0008f6a; 
			12'd544  : q <= 28'h0009874; 
			12'd545  : q <= 28'h0004c84; 
			12'd546  : q <= 28'h0888438; 
			12'd547  : q <= 28'hfd62f81; 
			12'd548  : q <= 28'h01c851e; 
			12'd549  : q <= 28'h00275ae; 
			12'd550  : q <= 28'hfff4e85; 
			12'd551  : q <= 28'hfe43582; 
			12'd552  : q <= 28'hffe937a; 
			12'd553  : q <= 28'h0018128; 
			12'd554  : q <= 28'h00e7fb9; 
			12'd555  : q <= 28'hffe3882; 
			12'd556  : q <= 28'h0017aad; 
			12'd557  : q <= 28'hff03182; 
			12'd558  : q <= 28'hffe997b; 
			12'd559  : q <= 28'h0005586; 
			12'd560  : q <= 28'hffda97d; 
			12'd561  : q <= 28'h000729b; 
			12'd562  : q <= 28'h0038a54; 
			12'd563  : q <= 28'hffbae75; 
			12'd564  : q <= 28'h0077693; 
			12'd565  : q <= 28'h0008443; 
			12'd566  : q <= 28'hff74087; 
			12'd567  : q <= 28'h000668d; 
			12'd568  : q <= 28'h0014aa2; 
			12'd569  : q <= 28'h0009f59; 
			12'd570  : q <= 28'h000398e; 
			12'd571  : q <= 28'h0005f97; 
			12'd572  : q <= 28'h0009055; 
			12'd573  : q <= 28'h0004e8d; 
			12'd574  : q <= 28'h000935e; 
			12'd575  : q <= 28'h000438b; 
			12'd576  : q <= 28'h002812d; 
			12'd577  : q <= 28'h0009571; 
			12'd578  : q <= 28'hfff4f88; 
			12'd579  : q <= 28'hffb5388; 
			12'd580  : q <= 28'hffdbc75; 
			12'd581  : q <= 28'h004863a; 
			12'd582  : q <= 28'h0008d61; 
			12'd583  : q <= 28'h0008a41; 
			12'd584  : q <= 28'h0008957; 
			12'd585  : q <= 28'hfff4d8a; 
			12'd586  : q <= 28'h0006690; 
			12'd587  : q <= 28'h0008e64; 
			12'd588  : q <= 28'h00d76b6; 
			12'd589  : q <= 28'hffc3b88; 
			12'd590  : q <= 28'hfff3b83; 
			12'd591  : q <= 28'h00077a5; 
			12'd592  : q <= 28'h001833c; 
			12'd593  : q <= 28'h0009f72; 
			12'd594  : q <= 28'hfff2f82; 
			12'd595  : q <= 28'h0258327; 
			12'd596  : q <= 28'h000885c; 
			12'd597  : q <= 28'h0009f7c; 
			12'd598  : q <= 28'h0006e95; 
			12'd599  : q <= 28'h0098624; 
			12'd600  : q <= 28'hfff5987; 
			12'd601  : q <= 28'h0007b9c; 
			12'd602  : q <= 28'hffa1d81; 
			12'd603  : q <= 28'h000a27a; 
			12'd604  : q <= 28'h000833f; 
			12'd605  : q <= 28'h0008a5e; 
			12'd606  : q <= 28'hff63082; 
			12'd607  : q <= 28'h000a57a; 
			12'd608  : q <= 28'h0009f73; 
			12'd609  : q <= 28'h0005f8a; 
			12'd610  : q <= 28'h02c801f; 
			12'd611  : q <= 28'h0005289; 
			12'd612  : q <= 28'h0006a92; 
			12'd613  : q <= 28'h000628e; 
			12'd614  : q <= 28'hffe3882; 
			12'd615  : q <= 28'h0008f6e; 
			12'd616  : q <= 28'h00776b2; 
			12'd617  : q <= 28'h002863a; 
			12'd618  : q <= 28'hfffa274; 
			12'd619  : q <= 28'h0018746; 
			12'd620  : q <= 28'hffa3481; 
			12'd621  : q <= 28'h000759c; 
			12'd622  : q <= 28'h0008133; 
			12'd623  : q <= 28'h0007b8b; 
			12'd624  : q <= 28'h00076ad; 
			12'd625  : q <= 28'h0008957; 
			12'd626  : q <= 28'hffb0680; 
			12'd627  : q <= 28'h0038528; 
			12'd628  : q <= 28'hffeba76; 
			12'd629  : q <= 28'h0028e64; 
			12'd630  : q <= 28'hfffae76; 
			12'd631  : q <= 28'hff24185; 
			12'd632  : q <= 28'h002844e; 
			12'd633  : q <= 28'hffd2184; 
			12'd634  : q <= 28'h000926c; 
			12'd635  : q <= 28'h0008768; 
			12'd636  : q <= 28'h000a875; 
			12'd637  : q <= 28'h0005c84; 
			12'd638  : q <= 28'hffd2081; 
			12'd639  : q <= 28'h000a179; 
			12'd640  : q <= 28'hfc82681; 
			12'd641  : q <= 28'h0016c91; 
			12'd642  : q <= 28'h000668f; 
			12'd643  : q <= 28'hfff997b; 
			12'd644  : q <= 28'h0005987; 
			12'd645  : q <= 28'h0017697; 
			12'd646  : q <= 28'h01f8011; 
			12'd647  : q <= 28'hffd967e; 
			12'd648  : q <= 28'h0016f96; 
			12'd649  : q <= 28'h0006e8a; 
			12'd650  : q <= 28'hffc3081; 
			12'd651  : q <= 28'h000876c; 
			12'd652  : q <= 28'hfffa274; 
			12'd653  : q <= 28'h001844d; 
			12'd654  : q <= 28'h0018241; 
			12'd655  : q <= 28'h0007896; 
			12'd656  : q <= 28'h0028127; 
			12'd657  : q <= 28'hfffa67d; 
			12'd658  : q <= 28'h0009f73; 
			12'd659  : q <= 28'hffe578a; 
			12'd660  : q <= 28'hff73081; 
			12'd661  : q <= 28'h000618a; 
			12'd662  : q <= 28'hff3af75; 
			12'd663  : q <= 28'h0018c73; 
			12'd664  : q <= 28'hfff5687; 
			12'd665  : q <= 28'h000a679; 
			12'd666  : q <= 28'h000678b; 
			12'd667  : q <= 28'hfffa37b; 
			12'd668  : q <= 28'hfff4c84; 
			12'd669  : q <= 28'h00780b7; 
			12'd670  : q <= 28'hffea676; 
			12'd671  : q <= 28'h00a833e; 
			12'd672  : q <= 28'h00275a3; 
			12'd673  : q <= 28'h000628c; 
			12'd674  : q <= 28'h0008345; 
			12'd675  : q <= 28'h0006789; 
			12'd676  : q <= 28'h003875f; 
			12'd677  : q <= 28'h0007ab0; 
			12'd678  : q <= 28'h0008964; 
			12'd679  : q <= 28'h00465b6; 
			12'd680  : q <= 28'h005569b; 
			12'd681  : q <= 28'h0005999; 
			12'd682  : q <= 28'h0025391; 
			12'd683  : q <= 28'h0004d8d; 
			12'd684  : q <= 28'h0005d91; 
			12'd685  : q <= 28'h0005489; 
			12'd686  : q <= 28'hfff458c; 
			12'd687  : q <= 28'h0028646; 
			12'd688  : q <= 28'hfef4a86; 
			12'd689  : q <= 28'h0009668; 
			12'd690  : q <= 28'h0005a8a; 
			12'd691  : q <= 28'h0008a59; 
			12'd692  : q <= 28'h00c8457; 
			12'd693  : q <= 28'h0005088; 
			12'd694  : q <= 28'h000718d; 
			12'd695  : q <= 28'h0004d86; 
			12'd696  : q <= 28'h0007aa9; 
			12'd697  : q <= 28'h0005187; 
			12'd698  : q <= 28'hfffa479; 
			12'd699  : q <= 28'hfff2682; 
			12'd700  : q <= 28'h0006e96; 
			12'd701  : q <= 28'h00479e8; 
			12'd702  : q <= 28'h0005a8e; 
			12'd703  : q <= 28'h00073a8; 
			12'd704  : q <= 28'h0009065; 
			12'd705  : q <= 28'h000895c; 
			12'd706  : q <= 28'h002862d; 
			12'd707  : q <= 28'hfff3a82; 
			12'd708  : q <= 28'h00076a9; 
			12'd709  : q <= 28'h000a171; 
			12'd710  : q <= 28'h0008a67; 
			12'd711  : q <= 28'h0018953; 
			12'd712  : q <= 28'hffdc77f; 
			12'd713  : q <= 28'h000875b; 
			12'd714  : q <= 28'h0007794; 
			12'd715  : q <= 28'h0008758; 
			12'd716  : q <= 28'h0037bbf; 
			12'd717  : q <= 28'h00073a3; 
			12'd718  : q <= 28'h001885b; 
			12'd719  : q <= 28'h0006c93; 
			12'd720  : q <= 28'hfff4c87; 
			12'd721  : q <= 28'h004812a; 
			12'd722  : q <= 28'h0017ab5; 
			12'd723  : q <= 28'h0018337; 
			12'd724  : q <= 28'hffd3186; 
			12'd725  : q <= 28'h000916b; 
			12'd726  : q <= 28'h0006c8b; 
			12'd727  : q <= 28'h0028240; 
			12'd728  : q <= 28'hff7b87c; 
			12'd729  : q <= 28'h000628a; 
			12'd730  : q <= 28'h0009774; 
			12'd731  : q <= 28'h0028347; 
			12'd732  : q <= 28'hffe9b76; 
			12'd733  : q <= 28'hfff5886; 
			12'd734  : q <= 28'h0009168; 
			12'd735  : q <= 28'h0006f94; 
			12'd736  : q <= 28'hfff2584; 
			12'd737  : q <= 28'h0008758; 
			12'd738  : q <= 28'h0007798; 
			12'd739  : q <= 28'h00177b3; 
			12'd740  : q <= 28'h0008c60; 
			12'd741  : q <= 28'hffc648b; 
			12'd742  : q <= 28'hff52983; 
			12'd743  : q <= 28'h0008347; 
			12'd744  : q <= 28'hfffa679; 
			12'd745  : q <= 28'hfff8d68; 
			12'd746  : q <= 28'h0005187; 
			12'd747  : q <= 28'hfffaf77; 
			12'd748  : q <= 28'h0008c73; 
			12'd749  : q <= 28'hffda375; 
			12'd750  : q <= 28'hffc4684; 
			12'd751  : q <= 28'hfff5584; 
			12'd752  : q <= 28'hffe987c; 
			12'd753  : q <= 28'h0006a8d; 
			12'd754  : q <= 28'h0028b6b; 
			12'd755  : q <= 28'hfffa474; 
			12'd756  : q <= 28'h0018539; 
			12'd757  : q <= 28'h0005084; 
			12'd758  : q <= 28'h0037cab; 
			12'd759  : q <= 28'h0005b86; 
			12'd760  : q <= 28'hffbe17f; 
			12'd761  : q <= 28'hfe82581; 
			12'd762  : q <= 28'h0018a6c; 
			12'd763  : q <= 28'h0006a8c; 
			12'd764  : q <= 28'h0037891; 
			12'd765  : q <= 28'hfffa072; 
			12'd766  : q <= 28'hfee4f85; 
			12'd767  : q <= 28'hfea1480; 
			12'd768  : q <= 28'h0078320; 
			12'd769  : q <= 28'h00b78bc; 
			12'd770  : q <= 28'hffd648d; 
			12'd771  : q <= 28'h003865e; 
			12'd772  : q <= 28'h000a278; 
			12'd773  : q <= 28'h0008860; 
			12'd774  : q <= 28'hfe42d85; 
			12'd775  : q <= 28'h0008862; 
			12'd776  : q <= 28'h0007693; 
			12'd777  : q <= 28'h0005284; 
			12'd778  : q <= 28'h0007aa5; 
			12'd779  : q <= 28'h0007099; 
			12'd780  : q <= 28'h000678c; 
			12'd781  : q <= 28'hff4a85f; 
			12'd782  : q <= 28'h0009458; 
			12'd783  : q <= 28'h0015c97; 
			12'd784  : q <= 28'h0008c49; 
			12'd785  : q <= 28'h000448b; 
			12'd786  : q <= 28'h0006292; 
			12'd787  : q <= 28'h0008c58; 
			12'd788  : q <= 28'h000548a; 
			12'd789  : q <= 28'h0005b89; 
			12'd790  : q <= 28'h0006d91; 
			12'd791  : q <= 28'h0008756; 
			12'd792  : q <= 28'h00074a0; 
			12'd793  : q <= 28'hffd3c83; 
			12'd794  : q <= 28'h000886a; 
			12'd795  : q <= 28'h0006d94; 
			12'd796  : q <= 28'hfff4a85; 
			12'd797  : q <= 28'h000875b; 
			12'd798  : q <= 28'h0017898; 
			12'd799  : q <= 28'hfff3682; 
			12'd800  : q <= 28'h0017aaf; 
			12'd801  : q <= 28'h002895f; 
			12'd802  : q <= 28'h0009262; 
			12'd803  : q <= 28'hfff5e88; 
			12'd804  : q <= 28'h0067f9b; 
			12'd805  : q <= 28'h0007199; 
			12'd806  : q <= 28'h002862f; 
			12'd807  : q <= 28'h0009b70; 
			12'd808  : q <= 28'hfff638f; 
			12'd809  : q <= 28'h0028134; 
			12'd810  : q <= 28'h000966b; 
			12'd811  : q <= 28'h0008d66; 
			12'd812  : q <= 28'h001548b; 
			12'd813  : q <= 28'h0008b64; 
			12'd814  : q <= 28'h0018f6b; 
			12'd815  : q <= 28'hfffab75; 
			12'd816  : q <= 28'h002894a; 
			12'd817  : q <= 28'h00377bb; 
			12'd818  : q <= 28'h000648a; 
			12'd819  : q <= 28'h0006c8f; 
			12'd820  : q <= 28'hffd5c87; 
			12'd821  : q <= 28'hfffaf76; 
			12'd822  : q <= 28'h000648a; 
			12'd823  : q <= 28'hffc3280; 
			12'd824  : q <= 28'h000688f; 
			12'd825  : q <= 28'h0007297; 
			12'd826  : q <= 28'h001885f; 
			12'd827  : q <= 28'h000824c; 
			12'd828  : q <= 28'hfff8d7b; 
			12'd829  : q <= 28'h00375a4; 
			12'd830  : q <= 28'h0088a57; 
			12'd831  : q <= 28'h0002b80; 
			12'd832  : q <= 28'h0008778; 
			12'd833  : q <= 28'h00176a4; 
			12'd834  : q <= 28'h0007b9a; 
			12'd835  : q <= 28'h0018452; 
			12'd836  : q <= 28'hffb6885; 
			12'd837  : q <= 28'h0008861; 
			12'd838  : q <= 28'h0009078; 
			12'd839  : q <= 28'h00074a0; 
			12'd840  : q <= 28'h0008854; 
			12'd841  : q <= 28'hfff1c80; 
			12'd842  : q <= 28'h000906e; 
			12'd843  : q <= 28'h0006a8b; 
			12'd844  : q <= 28'h0017cad; 
			12'd845  : q <= 28'h001865c; 
			12'd846  : q <= 28'h0038853; 
			12'd847  : q <= 28'h00176aa; 
			12'd848  : q <= 28'h0028c63; 
			12'd849  : q <= 28'h00078ba; 
			12'd850  : q <= 28'h000628b; 
			12'd851  : q <= 28'h0004182; 
			12'd852  : q <= 28'hffea57e; 
			12'd853  : q <= 28'h00d79c9; 
			12'd854  : q <= 28'h0008746; 
			12'd855  : q <= 28'h0008a67; 
			12'd856  : q <= 28'hffe9d7b; 
			12'd857  : q <= 28'h00178b3; 
			12'd858  : q <= 28'hfff4887; 
			12'd859  : q <= 28'h000b478; 
			12'd860  : q <= 28'h000638e; 
			12'd861  : q <= 28'h0005e86; 
			12'd862  : q <= 28'h0006289; 
			12'd863  : q <= 28'h00179be; 
			12'd864  : q <= 28'h0017b8f; 
			12'd865  : q <= 28'hffcb077; 
			12'd866  : q <= 28'h0008954; 
			12'd867  : q <= 28'h0078354; 
			12'd868  : q <= 28'h000779b; 
			12'd869  : q <= 28'h0007096; 
			12'd870  : q <= 28'h0008b6b; 
			12'd871  : q <= 28'h0008966; 
			12'd872  : q <= 28'h000906d; 
			12'd873  : q <= 28'h0008455; 
			12'd874  : q <= 28'h0407cb6; 
			12'd875  : q <= 28'hfff4582; 
			12'd876  : q <= 28'hff6af80; 
			12'd877  : q <= 28'h0006d8d; 
			12'd878  : q <= 28'h0006c89; 
			12'd879  : q <= 28'h00679c0; 
			12'd880  : q <= 28'hffe6c8d; 
			12'd881  : q <= 28'h0009873; 
			12'd882  : q <= 28'hfff698c; 
			12'd883  : q <= 28'h0017294; 
			12'd884  : q <= 28'h0008f71; 
			12'd885  : q <= 28'h00076a2; 
			12'd886  : q <= 28'h0007497; 
			12'd887  : q <= 28'h0008863; 
			12'd888  : q <= 28'h0008a5f; 
			12'd889  : q <= 28'h0006e8f; 
			12'd890  : q <= 28'hffb2d84; 
			12'd891  : q <= 28'h0006f91; 
			12'd892  : q <= 28'h005843c; 
			12'd893  : q <= 28'h0009972; 
			12'd894  : q <= 28'hffe6986; 
			12'd895  : q <= 28'h0008456; 
			12'd896  : q <= 28'hffeb07c; 
			12'd897  : q <= 28'h0008458; 
			12'd898  : q <= 28'hffd2a84; 
			12'd899  : q <= 28'h0006f90; 
			12'd900  : q <= 28'hff8c77e; 
			12'd901  : q <= 28'hffd2880; 
			12'd902  : q <= 28'h0228446; 
			12'd903  : q <= 28'h0005f85; 
			12'd904  : q <= 28'h0009573; 
			12'd905  : q <= 28'h00779bb; 
			12'd906  : q <= 28'h0008769; 
			12'd907  : q <= 28'h0137f20; 
			12'd908  : q <= 28'hffc0d84; 
			12'd909  : q <= 28'hfffae77; 
			12'd910  : q <= 28'h000997a; 
			12'd911  : q <= 28'h0005685; 
			12'd912  : q <= 28'hfff6f86; 
			12'd913  : q <= 28'h008813e; 
			12'd914  : q <= 28'h0009279; 
			12'd915  : q <= 28'hff96386; 
			12'd916  : q <= 28'h00b539f; 
			12'd917  : q <= 28'h0026cb1; 
			12'd918  : q <= 28'h0005f97; 
			12'd919  : q <= 28'h0003487; 
			12'd920  : q <= 28'h0008a4f; 
			12'd921  : q <= 28'h0008758; 
			12'd922  : q <= 28'h0008754; 
			12'd923  : q <= 28'h0009362; 
			12'd924  : q <= 28'h0006e9d; 
			12'd925  : q <= 28'hfff4b88; 
			12'd926  : q <= 28'h0008c62; 
			12'd927  : q <= 28'h0006d93; 
			12'd928  : q <= 28'h0005f8c; 
			12'd929  : q <= 28'h000749c; 
			12'd930  : q <= 28'h0004c84; 
			12'd931  : q <= 28'hfffab78; 
			12'd932  : q <= 28'h0005686; 
			12'd933  : q <= 28'h0018a64; 
			12'd934  : q <= 28'h000729c; 
			12'd935  : q <= 28'h0005f88; 
			12'd936  : q <= 28'hfff9a72; 
			12'd937  : q <= 28'hffd4888; 
			12'd938  : q <= 28'h0008556; 
			12'd939  : q <= 28'h0158314; 
			12'd940  : q <= 28'h0005484; 
			12'd941  : q <= 28'h002863b; 
			12'd942  : q <= 28'h000936d; 
			12'd943  : q <= 28'h0006f8e; 
			12'd944  : q <= 28'h00775a8; 
			12'd945  : q <= 28'h002875e; 
			12'd946  : q <= 28'hffeb576; 
			12'd947  : q <= 28'h0018745; 
			12'd948  : q <= 28'h001813e; 
			12'd949  : q <= 28'h0006d8e; 
			12'd950  : q <= 28'h0008d69; 
			12'd951  : q <= 28'hffaaf7c; 
			12'd952  : q <= 28'h0005f87; 
			12'd953  : q <= 28'h0009b76; 
			12'd954  : q <= 28'h004812e; 
			12'd955  : q <= 28'hfff2985; 
			12'd956  : q <= 28'h000729e; 
			12'd957  : q <= 28'h0008c6e; 
			12'd958  : q <= 28'hffe1d80; 
			12'd959  : q <= 28'h0017aac; 
			12'd960  : q <= 28'h0005884; 
			12'd961  : q <= 28'h0007a9f; 
			12'd962  : q <= 28'hfff9470; 
			12'd963  : q <= 28'h000638b; 
			12'd964  : q <= 28'hffe2a7f; 
			12'd965  : q <= 28'hffe6887; 
			12'd966  : q <= 28'h0009e75; 
			12'd967  : q <= 28'h0018e6a; 
			12'd968  : q <= 28'h000906f; 
			12'd969  : q <= 28'h0007bac; 
			12'd970  : q <= 28'h0088130; 
			12'd971  : q <= 28'hfec3c86; 
			12'd972  : q <= 28'h0018147; 
			12'd973  : q <= 28'h0009f78; 
			12'd974  : q <= 28'h0005484; 
			12'd975  : q <= 28'hfe43c84; 
			12'd976  : q <= 28'h0006889; 
			12'd977  : q <= 28'h0008c6f; 
			12'd978  : q <= 28'h0008d6b; 
			12'd979  : q <= 28'h0008b79; 
			12'd980  : q <= 28'h0018457; 
			12'd981  : q <= 28'h00080a2; 
			12'd982  : q <= 28'h0008d6c; 
			12'd983  : q <= 28'hfff718b; 
			12'd984  : q <= 28'h000b678; 
			12'd985  : q <= 28'h000688a; 
			12'd986  : q <= 28'hffac979; 
			12'd987  : q <= 28'h0006d8e; 
			12'd988  : q <= 28'h00178b3; 
			12'd989  : q <= 28'h0068661; 
			12'd990  : q <= 28'h009802b; 
			12'd991  : q <= 28'h0027ba3; 
			12'd992  : q <= 28'h0009772; 
			12'd993  : q <= 28'h001864c; 
			12'd994  : q <= 28'h0004d82; 
			12'd995  : q <= 28'h0006986; 
			12'd996  : q <= 28'hffe9473; 
			12'd997  : q <= 28'h0028644; 
			12'd998  : q <= 28'h00777b5; 
			12'd999  : q <= 28'h0018a60; 
			12'd1000 : q <= 28'hffa6086; 
			12'd1001 : q <= 28'h0006e94; 
			12'd1002 : q <= 28'h0008763; 
			12'd1003 : q <= 28'h0027d91; 
			12'd1004 : q <= 28'h0008e6e; 
			12'd1005 : q <= 28'h000906f; 
			12'd1006 : q <= 28'h0009b74; 
			12'd1007 : q <= 28'h0008969; 
			12'd1008 : q <= 28'h0006f92; 
			12'd1009 : q <= 28'hffc4d85; 
			12'd1010 : q <= 28'h0008761; 
			12'd1011 : q <= 28'h000886c; 
			12'd1012 : q <= 28'h0008c6b; 
			12'd1013 : q <= 28'hfe32485; 
			12'd1014 : q <= 28'hffdc678; 
			12'd1015 : q <= 28'h0008954; 
			12'd1016 : q <= 28'h0009372; 
			12'd1017 : q <= 28'h001855d; 
			12'd1018 : q <= 28'h0057f28; 
			12'd1019 : q <= 28'h00079a0; 
			12'd1020 : q <= 28'h0008864; 
			12'd1021 : q <= 28'hfffac80; 
			12'd1022 : q <= 28'hfff4f83; 
			12'd1023 : q <= 28'h0007d93; 
			12'd1024 : q <= 28'h0009a74; 
			12'd1025 : q <= 28'h0118637; 
			12'd1026 : q <= 28'h0068035; 
			12'd1027 : q <= 28'h0007cb5; 
			12'd1028 : q <= 28'h0005783; 
			12'd1029 : q <= 28'h0008e71; 
			12'd1030 : q <= 28'hffea376; 
			12'd1031 : q <= 28'h000608b; 
			12'd1032 : q <= 28'hfff5483; 
			12'd1033 : q <= 28'h0007da4; 
			12'd1034 : q <= 28'hfe72780; 
			12'd1035 : q <= 28'hfa70f84; 
			12'd1036 : q <= 28'hff5b277; 
			12'd1037 : q <= 28'h012841a; 
			12'd1038 : q <= 28'h0006d8d; 
			12'd1039 : q <= 28'h0007687; 
			12'd1040 : q <= 28'h0008764; 
			12'd1041 : q <= 28'h0009079; 
			12'd1042 : q <= 28'h0006e8d; 
			12'd1043 : q <= 28'hfff2484; 
			12'd1044 : q <= 28'h000708f; 
			12'd1045 : q <= 28'h0008878; 
			12'd1046 : q <= 28'h0008561; 
			12'd1047 : q <= 28'h0007a9c; 
			12'd1048 : q <= 28'h0006c8a; 
			12'd1049 : q <= 28'h0008b6b; 
			12'd1050 : q <= 28'h0009372; 
			12'd1051 : q <= 28'hffda378; 
			12'd1052 : q <= 28'h0008865; 
			12'd1053 : q <= 28'hffaa763; 
			12'd1054 : q <= 28'h0015f98; 
			12'd1055 : q <= 28'h0018a41; 
			12'd1056 : q <= 28'h0003f89; 
			12'd1057 : q <= 28'h0008f5a; 
			12'd1058 : q <= 28'h0006593; 
			12'd1059 : q <= 28'h0005e8d; 
			12'd1060 : q <= 28'hfff5f8e; 
			12'd1061 : q <= 28'hffbbf75; 
			12'd1062 : q <= 28'h0009063; 
			12'd1063 : q <= 28'h0005686; 
			12'd1064 : q <= 28'h0008d5f; 
			12'd1065 : q <= 28'h0008f69; 
			12'd1066 : q <= 28'h0005b88; 
			12'd1067 : q <= 28'h0008a60; 
			12'd1068 : q <= 28'hffba278; 
			12'd1069 : q <= 28'h000648e; 
			12'd1070 : q <= 28'hffe4185; 
			12'd1071 : q <= 28'h000844e; 
			12'd1072 : q <= 28'h0028949; 
			12'd1073 : q <= 28'h0006f95; 
			12'd1074 : q <= 28'h0038749; 
			12'd1075 : q <= 28'hffdb376; 
			12'd1076 : q <= 28'hffc4c86; 
			12'd1077 : q <= 28'h0006e97; 
			12'd1078 : q <= 28'h0028750; 
			12'd1079 : q <= 28'hffd4482; 
			12'd1080 : q <= 28'h0008b5f; 
			12'd1081 : q <= 28'h00178be; 
			12'd1082 : q <= 28'hfff3487; 
			12'd1083 : q <= 28'h0018459; 
			12'd1084 : q <= 28'hffeae7e; 
			12'd1085 : q <= 28'h0148139; 
			12'd1086 : q <= 28'hfda4b86; 
			12'd1087 : q <= 28'h00077b5; 
			12'd1088 : q <= 28'h0007a91; 
			12'd1089 : q <= 28'h0006d92; 
			12'd1090 : q <= 28'h001874f; 
			12'd1091 : q <= 28'h0005e86; 
			12'd1092 : q <= 28'hfe03c86; 
			12'd1093 : q <= 28'hfffb678; 
			12'd1094 : q <= 28'hffe728a; 
			12'd1095 : q <= 28'h0009871; 
			12'd1096 : q <= 28'h0008965; 
			12'd1097 : q <= 28'h0006086; 
			12'd1098 : q <= 28'h000a179; 
			12'd1099 : q <= 28'h0008556; 
			12'd1100 : q <= 28'h08b841e; 
			12'd1101 : q <= 28'h0047f23; 
			12'd1102 : q <= 28'hffdb67d; 
			12'd1103 : q <= 28'hfff3a81; 
			12'd1104 : q <= 28'h000769a; 
			12'd1105 : q <= 28'hfffa575; 
			12'd1106 : q <= 28'hffa2585; 
			12'd1107 : q <= 28'h0008356; 
			12'd1108 : q <= 28'hffe4687; 
			12'd1109 : q <= 28'h0008865; 
			12'd1110 : q <= 28'h0008968; 
			12'd1111 : q <= 28'h00177b0; 
			12'd1112 : q <= 28'h0008b5c; 
			12'd1113 : q <= 28'hfec2a80; 
			12'd1114 : q <= 28'h0058333; 
			12'd1115 : q <= 28'h00176a2; 
			12'd1116 : q <= 28'hfff977c; 
			12'd1117 : q <= 28'h0006388; 
			12'd1118 : q <= 28'h0006a8f; 
			12'd1119 : q <= 28'h0004f83; 
			12'd1120 : q <= 28'hfff6585; 
			12'd1121 : q <= 28'hffea075; 
			12'd1122 : q <= 28'hffc3586; 
			12'd1123 : q <= 28'h0008560; 
			12'd1124 : q <= 28'h0009476; 
			12'd1125 : q <= 28'h0007095; 
			12'd1126 : q <= 28'h000886b; 
			12'd1127 : q <= 28'h0005f86; 
			12'd1128 : q <= 28'h0007689; 
			12'd1129 : q <= 28'h001813c; 
			12'd1130 : q <= 28'hffcba81; 
			12'd1131 : q <= 28'hffaaa77; 
			12'd1132 : q <= 28'h0007088; 
			12'd1133 : q <= 28'h0026f91; 
			12'd1134 : q <= 28'h0007287; 
			12'd1135 : q <= 28'h00279bf; 
			12'd1136 : q <= 28'h0008979; 
			12'd1137 : q <= 28'hffe2c80; 
			12'd1138 : q <= 28'hfffba7d; 
			12'd1139 : q <= 28'h0006688; 
			12'd1140 : q <= 28'h0008f7a; 
			12'd1141 : q <= 28'h00279c3; 
			12'd1142 : q <= 28'h0028a6b; 
			12'd1143 : q <= 28'h0006c8a; 
			12'd1144 : q <= 28'h0006c8a; 
			12'd1145 : q <= 28'hffd9674; 
			12'd1146 : q <= 28'hffa4384; 
			12'd1147 : q <= 28'h000bc79; 
			12'd1148 : q <= 28'hffd4684; 
			12'd1149 : q <= 28'h0005983; 
			12'd1150 : q <= 28'h0009077; 
			12'd1151 : q <= 28'h005769d; 
			12'd1152 : q <= 28'hfe84c84; 
			12'd1153 : q <= 28'h001814d; 
			12'd1154 : q <= 28'h0017cb0; 
			12'd1155 : q <= 28'hffe2a80; 
			12'd1156 : q <= 28'hfff4486; 
			12'd1157 : q <= 28'hffeb779; 
			12'd1158 : q <= 28'h002853d; 
			12'd1159 : q <= 28'h0009271; 
			12'd1160 : q <= 28'h0018c6a; 
			12'd1161 : q <= 28'h0277f0f; 
			12'd1162 : q <= 28'h000788a; 
			12'd1163 : q <= 28'h0006887; 
			12'd1164 : q <= 28'hffe9c7e; 
			12'd1165 : q <= 28'h00b8149; 
			12'd1166 : q <= 28'h0007ca1; 
			12'd1167 : q <= 28'hfe20f7f; 
			12'd1168 : q <= 28'h0008978; 
			12'd1169 : q <= 28'hfcb0f7f; 
			12'd1170 : q <= 28'h0007889; 
			12'd1171 : q <= 28'h0006f8d; 
			12'd1172 : q <= 28'h000947b; 
			12'd1173 : q <= 28'h0008767; 
			12'd1174 : q <= 28'h0006086; 
			12'd1175 : q <= 28'h0027ac4; 
			12'd1176 : q <= 28'h003864e; 
			12'd1177 : q <= 28'hfcaac78; 
			12'd1178 : q <= 28'h0009070; 
			12'd1179 : q <= 28'h0007396; 
			12'd1180 : q <= 28'h0009b7e; 
			12'd1181 : q <= 28'h0009973; 
			12'd1182 : q <= 28'h0006b85; 
			12'd1183 : q <= 28'h006855b; 
			12'd1184 : q <= 28'h0005085; 
			12'd1185 : q <= 28'h0005683; 
			12'd1186 : q <= 28'hffc957d; 
			12'd1187 : q <= 28'hffd9d76; 
			12'd1188 : q <= 28'h008842b; 
			12'd1189 : q <= 28'h0005783; 
			12'd1190 : q <= 28'hffe9c7f; 
			12'd1191 : q <= 28'h0006e8e; 
			12'd1192 : q <= 28'h0027c8b; 
			12'd1193 : q <= 28'h0025598; 
			12'd1194 : q <= 28'h000598e; 
			12'd1195 : q <= 28'h0008d54; 
			12'd1196 : q <= 28'h0005c8d; 
			12'd1197 : q <= 28'h0005a8e; 
			12'd1198 : q <= 28'h0006490; 
			12'd1199 : q <= 28'h02477b3; 
			12'd1200 : q <= 28'hfff4e87; 
			12'd1201 : q <= 28'h0008f67; 
			12'd1202 : q <= 28'h000865b; 
			12'd1203 : q <= 28'hffdaa76; 
			12'd1204 : q <= 28'h0008d63; 
			12'd1205 : q <= 28'h0005c88; 
			12'd1206 : q <= 28'h0007689; 
			12'd1207 : q <= 28'h0018353; 
			12'd1208 : q <= 28'hffeab7a; 
			12'd1209 : q <= 28'h000678b; 
			12'd1210 : q <= 28'h000a57a; 
			12'd1211 : q <= 28'h000865a; 
			12'd1212 : q <= 28'hfff6189; 
			12'd1213 : q <= 28'h0008863; 
			12'd1214 : q <= 28'h0005b87; 
			12'd1215 : q <= 28'h00277af; 
			12'd1216 : q <= 28'h00a8311; 
			12'd1217 : q <= 28'h0004d83; 
			12'd1218 : q <= 28'hfffa47d; 
			12'd1219 : q <= 28'h0008761; 
			12'd1220 : q <= 28'h000778a; 
			12'd1221 : q <= 28'hfff4882; 
			12'd1222 : q <= 28'hffd4c83; 
			12'd1223 : q <= 28'h000906f; 
			12'd1224 : q <= 28'h0007089; 
			12'd1225 : q <= 28'h0005784; 
			12'd1226 : q <= 28'h002769c; 
			12'd1227 : q <= 28'hffe4881; 
			12'd1228 : q <= 28'h0068544; 
			12'd1229 : q <= 28'h00477ac; 
			12'd1230 : q <= 28'h0058538; 
			12'd1231 : q <= 28'h0009b74; 
			12'd1232 : q <= 28'hffe7686; 
			12'd1233 : q <= 28'h0028764; 
			12'd1234 : q <= 28'hfeec67f; 
			12'd1235 : q <= 28'hfff3e81; 
			12'd1236 : q <= 28'hffe927b; 
			12'd1237 : q <= 28'h00f8040; 
			12'd1238 : q <= 28'h0009b7d; 
			12'd1239 : q <= 28'h0018038; 
			12'd1240 : q <= 28'h000a97e; 
			12'd1241 : q <= 28'h00a845f; 
			12'd1242 : q <= 28'h0007894; 
			12'd1243 : q <= 28'h0006185; 
			12'd1244 : q <= 28'hffe4b85; 
			12'd1245 : q <= 28'hfffbc78; 
			12'd1246 : q <= 28'h0008b6c; 
			12'd1247 : q <= 28'h000708f; 
			12'd1248 : q <= 28'h000799d; 
			12'd1249 : q <= 28'h0009a73; 
			12'd1250 : q <= 28'h0003e87; 
			12'd1251 : q <= 28'h0005f86; 
			12'd1252 : q <= 28'h0008c68; 
			12'd1253 : q <= 28'hfff367f; 
			12'd1254 : q <= 28'h0007794; 
			12'd1255 : q <= 28'h000708e; 
			12'd1256 : q <= 28'h00c8652; 
			12'd1257 : q <= 28'hfff9b74; 
			12'd1258 : q <= 28'hffd3483; 
			12'd1259 : q <= 28'h000865f; 
			12'd1260 : q <= 28'h0077e98; 
			12'd1261 : q <= 28'h000886a; 
			12'd1262 : q <= 28'h000788d; 
			12'd1263 : q <= 28'hffdad77; 
			12'd1264 : q <= 28'hfff5c85; 
			12'd1265 : q <= 28'h000875d; 
			12'd1266 : q <= 28'h0268438; 
			12'd1267 : q <= 28'h0017093; 
			12'd1268 : q <= 28'h0028a60; 
			12'd1269 : q <= 28'h0006f8f; 
			12'd1270 : q <= 28'h0006c8d; 
			12'd1271 : q <= 28'h0007397; 
			12'd1272 : q <= 28'h00b8750; 
			12'd1273 : q <= 28'h0007295; 
			12'd1274 : q <= 28'hfff748c; 
			12'd1275 : q <= 28'h0008861; 
			12'd1276 : q <= 28'h0009175; 
			12'd1277 : q <= 28'h0007190; 
			12'd1278 : q <= 28'h0006d8a; 
			12'd1279 : q <= 28'hff4b078; 
			12'd1280 : q <= 28'hff73884; 
			12'd1281 : q <= 28'h0008359; 
			12'd1282 : q <= 28'h0007ba4; 
			12'd1283 : q <= 28'h0006486; 
			12'd1284 : q <= 28'h00382d7; 
			12'd1285 : q <= 28'h0008d6e; 
			12'd1286 : q <= 28'h0006489; 
			12'd1287 : q <= 28'hfffbc79; 
			12'd1288 : q <= 28'h0108454; 
			12'd1289 : q <= 28'h0005e84; 
			12'd1290 : q <= 28'h00380ab; 
			12'd1291 : q <= 28'hffbad78; 
			12'd1292 : q <= 28'h0018667; 
			12'd1293 : q <= 28'h00078ab; 
			12'd1294 : q <= 28'h0006e88; 
			12'd1295 : q <= 28'h0027f29; 
			12'd1296 : q <= 28'h0006d90; 
			12'd1297 : q <= 28'hfffad78; 
			12'd1298 : q <= 28'h0008874; 
			12'd1299 : q <= 28'hfff9070; 
			12'd1300 : q <= 28'h0005f89; 
			12'd1301 : q <= 28'h000845f; 
			12'd1302 : q <= 28'hff74b84; 
			12'd1303 : q <= 28'h0006f8d; 
			12'd1304 : q <= 28'hff85285; 
			12'd1305 : q <= 28'hffe9874; 
			12'd1306 : q <= 28'h000798c; 
			12'd1307 : q <= 28'h0006e8c; 
			12'd1308 : q <= 28'hffc2884; 
			12'd1309 : q <= 28'h0007393; 
			12'd1310 : q <= 28'h0006a8b; 
			12'd1311 : q <= 28'h0006787; 
			12'd1312 : q <= 28'h0017a9c; 
			12'd1313 : q <= 28'hfff5b84; 
			12'd1314 : q <= 28'h003788e; 
			12'd1315 : q <= 28'hfff4481; 
			12'd1316 : q <= 28'h0638340; 
			12'd1317 : q <= 28'h0006d8a; 
			12'd1318 : q <= 28'hffc6385; 
			12'd1319 : q <= 28'h0008a6c; 
			12'd1320 : q <= 28'h0007da9; 
			12'd1321 : q <= 28'h0008767; 
			12'd1322 : q <= 28'h0009a7a; 
			12'd1323 : q <= 28'hfff6889; 
			12'd1324 : q <= 28'h0007c93; 
			12'd1325 : q <= 28'h000845b; 
			12'd1326 : q <= 28'h0009179; 
			12'd1327 : q <= 28'h00079b5; 
			12'd1328 : q <= 28'h0018647; 
			12'd1329 : q <= 28'hfff4881; 
			12'd1330 : q <= 28'hffebd7e; 
			12'd1331 : q <= 28'h0018357; 
			12'd1332 : q <= 28'h0017ea8; 
			12'd1333 : q <= 28'hfff3e80; 
			12'd1334 : q <= 28'h0009778; 
			12'd1335 : q <= 28'h0005d84; 
			12'd1336 : q <= 28'h0009a7e; 
			12'd1337 : q <= 28'hfff9474; 
			12'd1338 : q <= 28'h0008559; 
			12'd1339 : q <= 28'hffb3c80; 
			12'd1340 : q <= 28'hff9a67d; 
			12'd1341 : q <= 28'h0037091; 
			12'd1342 : q <= 28'h0006f88; 
			12'd1343 : q <= 28'h0008c6e; 
			12'd1344 : q <= 28'hffd6885; 
			12'd1345 : q <= 28'hff80c7f; 
			12'd1346 : q <= 28'h00d7caa; 
			12'd1347 : q <= 28'h0028a6c; 
			12'd1348 : q <= 28'h0007a8e; 
			12'd1349 : q <= 28'h000bd7a; 
			12'd1350 : q <= 28'h0008751; 
			12'd1351 : q <= 28'h00079b4; 
			12'd1352 : q <= 28'h0006188; 
			12'd1353 : q <= 28'h00e66ae; 
			12'd1354 : q <= 28'h0005598; 
			12'd1355 : q <= 28'h0008e59; 
			12'd1356 : q <= 28'h0006d91; 
			12'd1357 : q <= 28'h000598b; 
			12'd1358 : q <= 28'h000678c; 
			12'd1359 : q <= 28'h000618a; 
			12'd1360 : q <= 28'h000438a; 
			12'd1361 : q <= 28'h000618a; 
			12'd1362 : q <= 28'h000718b; 
			12'd1363 : q <= 28'h0005f8a; 
			12'd1364 : q <= 28'h0238d72; 
			12'd1365 : q <= 28'h0006d93; 
			12'd1366 : q <= 28'h0006f91; 
			12'd1367 : q <= 28'h0005685; 
			12'd1368 : q <= 28'h0007499; 
			12'd1369 : q <= 28'h000834b; 
			12'd1370 : q <= 28'h0006489; 
			12'd1371 : q <= 28'h0005e85; 
			12'd1372 : q <= 28'hffeba7d; 
			12'd1373 : q <= 28'h0006f91; 
			12'd1374 : q <= 28'hfff4285; 
			12'd1375 : q <= 28'hffcb177; 
			12'd1376 : q <= 28'h0018954; 
			12'd1377 : q <= 28'hfff3480; 
			12'd1378 : q <= 28'hffdae7d; 
			12'd1379 : q <= 28'h0008763; 
			12'd1380 : q <= 28'hfff926f; 
			12'd1381 : q <= 28'h0004882; 
			12'd1382 : q <= 28'h0005686; 
			12'd1383 : q <= 28'h0008764; 
			12'd1384 : q <= 28'h0008b64; 
			12'd1385 : q <= 28'hff83781; 
			12'd1386 : q <= 28'h000a57c; 
			12'd1387 : q <= 28'h001769f; 
			12'd1388 : q <= 28'h0048533; 
			12'd1389 : q <= 28'h0006687; 
			12'd1390 : q <= 28'h0007a90; 
			12'd1391 : q <= 28'hfe83480; 
			12'd1392 : q <= 28'hffbc481; 
			12'd1393 : q <= 28'hffdbf79; 
			12'd1394 : q <= 28'h0018966; 
			12'd1395 : q <= 28'hffb127f; 
			12'd1396 : q <= 28'hfd64985; 
			12'd1397 : q <= 28'h0006b89; 
			12'd1398 : q <= 28'hffea07c; 
			12'd1399 : q <= 28'h000845d; 
			12'd1400 : q <= 28'h0009675; 
			12'd1401 : q <= 28'h0005b83; 
			12'd1402 : q <= 28'hfff9977; 
			12'd1403 : q <= 28'hff85583; 
			12'd1404 : q <= 28'h0008e70; 
			12'd1405 : q <= 28'h000769d; 
			12'd1406 : q <= 28'h000a77f; 
			12'd1407 : q <= 28'h0008663; 
			12'd1408 : q <= 28'h0007694; 
			12'd1409 : q <= 28'hffe4481; 
			12'd1410 : q <= 28'h0008b6e; 
			12'd1411 : q <= 28'h00177ab; 
			12'd1412 : q <= 28'h0008756; 
			12'd1413 : q <= 28'h0006888; 
			12'd1414 : q <= 28'hfed3285; 
			12'd1415 : q <= 28'h0008b6c; 
			12'd1416 : q <= 28'hfff6d89; 
			12'd1417 : q <= 28'hfe4b078; 
			12'd1418 : q <= 28'h000738e; 
			12'd1419 : q <= 28'h000896c; 
			12'd1420 : q <= 28'hffaa47f; 
			12'd1421 : q <= 28'h0087f29; 
			12'd1422 : q <= 28'h0008a6c; 
			12'd1423 : q <= 28'h001759a; 
			12'd1424 : q <= 28'h0008771; 
			12'd1425 : q <= 28'h00078aa; 
			12'd1426 : q <= 28'h000708d; 
			12'd1427 : q <= 28'h0018354; 
			12'd1428 : q <= 28'h0005084; 
			12'd1429 : q <= 28'h0006987; 
			12'd1430 : q <= 28'hffc9e7b; 
			12'd1431 : q <= 28'h0005d84; 
			12'd1432 : q <= 28'hffb5984; 
			12'd1433 : q <= 28'h000845e; 
			12'd1434 : q <= 28'h00480ce; 
			12'd1435 : q <= 28'hffea577; 
			12'd1436 : q <= 28'hffd5386; 
			12'd1437 : q <= 28'h0008462; 
			12'd1438 : q <= 28'h0017d9e; 
			12'd1439 : q <= 28'hfc12f7f; 
			12'd1440 : q <= 28'h003855c; 
			12'd1441 : q <= 28'h0007293; 
			12'd1442 : q <= 28'h0007b95; 
			12'd1443 : q <= 28'hffd4080; 
			12'd1444 : q <= 28'hfff997c; 
			12'd1445 : q <= 28'h000835d; 
			12'd1446 : q <= 28'hffca97f; 
			12'd1447 : q <= 28'h00276a0; 
			12'd1448 : q <= 28'hfff5c87; 
			12'd1449 : q <= 28'h000718e; 
			12'd1450 : q <= 28'h0018442; 
			12'd1451 : q <= 28'hfff4780; 
			12'd1452 : q <= 28'h0017f90; 
			12'd1453 : q <= 28'h000718e; 
			12'd1454 : q <= 28'hfbb0783; 
			12'd1455 : q <= 28'hffd9171; 
			12'd1456 : q <= 28'hffe6e8c; 
			12'd1457 : q <= 28'h0005e83; 
			12'd1458 : q <= 28'h0017b9c; 
			12'd1459 : q <= 28'h0008869; 
			12'd1460 : q <= 28'h0007ba0; 
			12'd1461 : q <= 28'h002855c; 
			12'd1462 : q <= 28'h0037fac; 
			12'd1463 : q <= 28'h0006787; 
			12'd1464 : q <= 28'h0007797; 
			12'd1465 : q <= 28'h000739b; 
			12'd1466 : q <= 28'hfea4784; 
			12'd1467 : q <= 28'h0008768; 
			12'd1468 : q <= 28'h0008b74; 
			12'd1469 : q <= 28'h001886b; 
			12'd1470 : q <= 28'h0007392; 
			12'd1471 : q <= 28'h0007596; 
			12'd1472 : q <= 28'h0008755; 
			12'd1473 : q <= 28'h0037e22; 
			12'd1474 : q <= 28'h0078200; 
			12'd1475 : q <= 28'h00179b3; 
			12'd1476 : q <= 28'h0028554; 
			12'd1477 : q <= 28'h0009474; 
			12'd1478 : q <= 28'h0038a69; 
			12'd1479 : q <= 28'h0006c8a; 
			12'd1480 : q <= 28'h0028658; 
			12'd1481 : q <= 28'h0009072; 
			12'd1482 : q <= 28'h001886f; 
			12'd1483 : q <= 28'h00778a8; 
			12'd1484 : q <= 28'hffb0083; 
			12'd1485 : q <= 28'hfea067e; 
			12'd1486 : q <= 28'hffd5083; 
			12'd1487 : q <= 28'h0028040; 
			12'd1488 : q <= 28'hfffa37e; 
			12'd1489 : q <= 28'h000835e; 
			12'd1490 : q <= 28'h0018d6f; 
			12'd1491 : q <= 28'h0009d75; 
			12'd1492 : q <= 28'hfff9e7d; 
			12'd1493 : q <= 28'hffc237f; 
			12'd1494 : q <= 28'h001788c; 
			12'd1495 : q <= 28'h0003c80; 
			12'd1496 : q <= 28'h0009578; 
			12'd1497 : q <= 28'hfdc167f; 
			12'd1498 : q <= 28'h01b832c; 
			12'd1499 : q <= 28'hff3bc7a; 
			12'd1500 : q <= 28'hfff6387; 
			12'd1501 : q <= 28'h0008566; 
			12'd1502 : q <= 28'h0027eb8; 
			12'd1503 : q <= 28'h000718d; 
			12'd1504 : q <= 28'h0008a6a; 
			12'd1505 : q <= 28'h0009574; 
			12'd1506 : q <= 28'h0007587; 
			12'd1507 : q <= 28'h0006186; 
			12'd1508 : q <= 28'hfff997e; 
			12'd1509 : q <= 28'h000728f; 
			12'd1510 : q <= 28'h0008b71; 
			12'd1511 : q <= 28'hfff6986; 
			12'd1512 : q <= 28'h000947f; 
			12'd1513 : q <= 28'hfedd67b; 
			12'd1514 : q <= 28'hff63d84; 
			12'd1515 : q <= 28'h0006f8a; 
			12'd1516 : q <= 28'h0008b7d; 
			12'd1517 : q <= 28'hffe9375; 
			12'd1518 : q <= 28'h0048457; 
			12'd1519 : q <= 28'hff83880; 
			12'd1520 : q <= 28'h00181a8; 
			12'd1521 : q <= 28'hffe377f; 
			12'd1522 : q <= 28'h000808c; 
			12'd1523 : q <= 28'h0006986; 
			12'd1524 : q <= 28'h0008a7f; 
			12'd1525 : q <= 28'h0007596; 
			12'd1526 : q <= 28'h0008778; 
			12'd1527 : q <= 28'h0008360; 
			12'd1528 : q <= 28'h0067b94; 
			12'd1529 : q <= 28'h0008665; 
			12'd1530 : q <= 28'h0015998; 
			12'd1531 : q <= 28'hffeae72; 
			12'd1532 : q <= 28'h0008e5b; 
			12'd1533 : q <= 28'h000894e; 
			12'd1534 : q <= 28'h0005d88; 
			12'd1535 : q <= 28'hfff498c; 
			12'd1536 : q <= 28'h0008658; 
			12'd1537 : q <= 28'h002799f; 
			12'd1538 : q <= 28'hff75587; 
			12'd1539 : q <= 28'h001845e; 
			12'd1540 : q <= 28'h0004b82; 
			12'd1541 : q <= 28'h0045e8b; 
			12'd1542 : q <= 28'hfff5c85; 
			12'd1543 : q <= 28'h0009678; 
			12'd1544 : q <= 28'h0005183; 
			12'd1545 : q <= 28'hfffa17b; 
			12'd1546 : q <= 28'hfff3280; 
			12'd1547 : q <= 28'h0027eaf; 
			12'd1548 : q <= 28'h0018455; 
			12'd1549 : q <= 28'hfe23b86; 
			12'd1550 : q <= 28'h00777ac; 
			12'd1551 : q <= 28'h0018545; 
			12'd1552 : q <= 28'h000824a; 
			12'd1553 : q <= 28'h0027da3; 
			12'd1554 : q <= 28'h001855d; 
			12'd1555 : q <= 28'h0009d79; 
			12'd1556 : q <= 28'hffd4380; 
			12'd1557 : q <= 28'hfe63a84; 
			12'd1558 : q <= 28'hffeb278; 
			12'd1559 : q <= 28'h0008b6d; 
			12'd1560 : q <= 28'hfff9b75; 
			12'd1561 : q <= 28'h0028654; 
			12'd1562 : q <= 28'h000896a; 
			12'd1563 : q <= 28'h0006d87; 
			12'd1564 : q <= 28'h0006185; 
			12'd1565 : q <= 28'h0018669; 
			12'd1566 : q <= 28'hff8317f; 
			12'd1567 : q <= 28'hffe997e; 
			12'd1568 : q <= 28'h0038034; 
			12'd1569 : q <= 28'h0007c92; 
			12'd1570 : q <= 28'h001802e; 
			12'd1571 : q <= 28'h0008d7d; 
			12'd1572 : q <= 28'hffd6a89; 
			12'd1573 : q <= 28'h0017f93; 
			12'd1574 : q <= 28'h0008868; 
			12'd1575 : q <= 28'hffd9381; 
			12'd1576 : q <= 28'h000759a; 
			12'd1577 : q <= 28'h000708a; 
			12'd1578 : q <= 28'h000845e; 
			12'd1579 : q <= 28'hffe9b7c; 
			12'd1580 : q <= 28'hfff5482; 
			12'd1581 : q <= 28'h0017b9c; 
			12'd1582 : q <= 28'h00277a7; 
			12'd1583 : q <= 28'h009852b; 
			12'd1584 : q <= 28'h001845f; 
			12'd1585 : q <= 28'hfffa47f; 
			12'd1586 : q <= 28'h0009672; 
			12'd1587 : q <= 28'h0008b58; 
			12'd1588 : q <= 28'hffe3680; 
			12'd1589 : q <= 28'h0008975; 
			12'd1590 : q <= 28'h0009373; 
			12'd1591 : q <= 28'h0008a6c; 
			12'd1592 : q <= 28'hffe6886; 
			12'd1593 : q <= 28'hfff6c8c; 
			12'd1594 : q <= 28'hff7a877; 
			12'd1595 : q <= 28'h0006c8e; 
			12'd1596 : q <= 28'h0008668; 
			12'd1597 : q <= 28'h0007796; 
			12'd1598 : q <= 28'h0009272; 
			12'd1599 : q <= 28'h001864a; 
			12'd1600 : q <= 28'h0006385; 
			12'd1601 : q <= 28'h000947e; 
			12'd1602 : q <= 28'hfff3c80; 
			12'd1603 : q <= 28'h0007c8f; 
			12'd1604 : q <= 28'h0008460; 
			12'd1605 : q <= 28'h0008b7c; 
			12'd1606 : q <= 28'h00078ab; 
			12'd1607 : q <= 28'h0148445; 
			12'd1608 : q <= 28'h0147f2d; 
			12'd1609 : q <= 28'h0028452; 
			12'd1610 : q <= 28'h0006787; 
			12'd1611 : q <= 28'hfff5884; 
			12'd1612 : q <= 28'h000759b; 
			12'd1613 : q <= 28'hffb2b85; 
			12'd1614 : q <= 28'h0006285; 
			12'd1615 : q <= 28'h0008d6f; 
			12'd1616 : q <= 28'hffbcc7a; 
			12'd1617 : q <= 28'h0006889; 
			12'd1618 : q <= 28'h0008c6f; 
			12'd1619 : q <= 28'h0007f95; 
			12'd1620 : q <= 28'h000ac78; 
			12'd1621 : q <= 28'h0008a6f; 
			12'd1622 : q <= 28'hfff397f; 
			12'd1623 : q <= 28'hffea07e; 
			12'd1624 : q <= 28'h0006586; 
			12'd1625 : q <= 28'h0047994; 
			12'd1626 : q <= 28'hffd9a74; 
			12'd1627 : q <= 28'h0006d8d; 
			12'd1628 : q <= 28'h0008560; 
			12'd1629 : q <= 28'hfffa37b; 
			12'd1630 : q <= 28'h001896a; 
			12'd1631 : q <= 28'h0007687; 
			12'd1632 : q <= 28'h00978a5; 
			12'd1633 : q <= 28'h0028538; 
			12'd1634 : q <= 28'hfd9297e; 
			12'd1635 : q <= 28'h0009378; 
			12'd1636 : q <= 28'h0006585; 
			12'd1637 : q <= 28'h0009a7b; 
			12'd1638 : q <= 28'h0006685; 
			12'd1639 : q <= 28'h0007893; 
			12'd1640 : q <= 28'h0006986; 
			12'd1641 : q <= 28'h005852d; 
			12'd1642 : q <= 28'hfffa878; 
			12'd1643 : q <= 28'h0068356; 
			12'd1644 : q <= 28'h000a878; 
			12'd1645 : q <= 28'h00e8347; 
			12'd1646 : q <= 28'h0006284; 
			12'd1647 : q <= 28'h004829e; 
			12'd1648 : q <= 28'h001835e; 
			12'd1649 : q <= 28'hfff997b; 
			12'd1650 : q <= 28'h0007392; 
			12'd1651 : q <= 28'h0005986; 
			12'd1652 : q <= 28'hffc1c7f; 
			12'd1653 : q <= 28'h0028370; 
			12'd1654 : q <= 28'h0006886; 
			12'd1655 : q <= 28'hff5a380; 
			12'd1656 : q <= 28'h00278ab; 
			12'd1657 : q <= 28'hfff7488; 
			12'd1658 : q <= 28'h0006e8b; 
			12'd1659 : q <= 28'h000758d; 
			12'd1660 : q <= 28'h0006e8a; 
			12'd1661 : q <= 28'h001865a; 
			12'd1662 : q <= 28'hffe9a76; 
			12'd1663 : q <= 28'h000758d; 
			12'd1664 : q <= 28'h0006988; 
			12'd1665 : q <= 28'h000678a; 
			12'd1666 : q <= 28'h0007390; 
			12'd1667 : q <= 28'h0028445; 
			12'd1668 : q <= 28'hfff327f; 
			12'd1669 : q <= 28'hfffaa80; 
			12'd1670 : q <= 28'hfff6384; 
			12'd1671 : q <= 28'h0007a90; 
			12'd1672 : q <= 28'h0008565; 
			12'd1673 : q <= 28'hff69d80; 
			12'd1674 : q <= 28'h0006585; 
			12'd1675 : q <= 28'h0007f98; 
			12'd1676 : q <= 28'h0027f29; 
			12'd1677 : q <= 28'h000977e; 
			12'd1678 : q <= 28'h0006b88; 
			12'd1679 : q <= 28'h0018a7d; 
			12'd1680 : q <= 28'h0005f83; 
			12'd1681 : q <= 28'hff6a581; 
			12'd1682 : q <= 28'h00077a3; 
			12'd1683 : q <= 28'h0008b6a; 
			12'd1684 : q <= 28'h0005e83; 
			12'd1685 : q <= 28'hffd9a7b; 
			12'd1686 : q <= 28'hfe7337f; 
			12'd1687 : q <= 28'hffc927d; 
			12'd1688 : q <= 28'h0006b8a; 
			12'd1689 : q <= 28'h0228360; 
			12'd1690 : q <= 28'hffab379; 
			12'd1691 : q <= 28'h0006e8a; 
			12'd1692 : q <= 28'h0009876; 
			12'd1693 : q <= 28'hfff9e7d; 
			12'd1694 : q <= 28'h0008666; 
			12'd1695 : q <= 28'h00b8644; 
			12'd1696 : q <= 28'hffb367f; 
			12'd1697 : q <= 28'h0007b8d; 
			12'd1698 : q <= 28'h000a578; 
			12'd1699 : q <= 28'hfff7587; 
			12'd1700 : q <= 28'h0008567; 
			12'd1701 : q <= 28'h0008e7a; 
			12'd1702 : q <= 28'h0008566; 
			12'd1703 : q <= 28'hff1a180; 
			12'd1704 : q <= 28'hfefb97a; 
			12'd1705 : q <= 28'hfee3a84; 
			12'd1706 : q <= 28'h0008668; 
			12'd1707 : q <= 28'h0007a8b; 
			12'd1708 : q <= 28'hffab67a; 
			12'd1709 : q <= 28'hffd4386; 
			12'd1710 : q <= 28'h0005c82; 
			12'd1711 : q <= 28'h000788b; 
			12'd1712 : q <= 28'h00362a4; 
			12'd1713 : q <= 28'h00670ac; 
			12'd1714 : q <= 28'h0008c57; 
			12'd1715 : q <= 28'h000528a; 
			12'd1716 : q <= 28'h001824b; 
			12'd1717 : q <= 28'h0006a88; 
			12'd1718 : q <= 28'h0004a83; 
			12'd1719 : q <= 28'h0006d8e; 
			12'd1720 : q <= 28'h000678a; 
			12'd1721 : q <= 28'h0006d8c; 
			12'd1722 : q <= 28'h0006589; 
			12'd1723 : q <= 28'h0007986; 
			12'd1724 : q <= 28'h0008f6c; 
			12'd1725 : q <= 28'h0008579; 
			12'd1726 : q <= 28'h000668b; 
			12'd1727 : q <= 28'h002779a; 
			12'd1728 : q <= 28'hffe5985; 
			12'd1729 : q <= 28'h0009e79; 
			12'd1730 : q <= 28'h0008762; 
			12'd1731 : q <= 28'h0008958; 
			12'd1732 : q <= 28'h000749e; 
			12'd1733 : q <= 28'h0005e88; 
			12'd1734 : q <= 28'h0006587; 
			12'd1735 : q <= 28'hff5b37f; 
			12'd1736 : q <= 28'h0088146; 
			12'd1737 : q <= 28'h0004487; 
			12'd1738 : q <= 28'h0007599; 
			12'd1739 : q <= 28'hffb5186; 
			12'd1740 : q <= 28'h0008667; 
			12'd1741 : q <= 28'h0008875; 
			12'd1742 : q <= 28'h001759a; 
			12'd1743 : q <= 28'hffd7189; 
			12'd1744 : q <= 28'h00177a4; 
			12'd1745 : q <= 28'h0005e88; 
			12'd1746 : q <= 28'h00378b6; 
			12'd1747 : q <= 28'h0007389; 
			12'd1748 : q <= 28'h000708d; 
			12'd1749 : q <= 28'h0007798; 
			12'd1750 : q <= 28'h000824d; 
			12'd1751 : q <= 28'h0008f72; 
			12'd1752 : q <= 28'hfff387f; 
			12'd1753 : q <= 28'hffca780; 
			12'd1754 : q <= 28'h0247f25; 
			12'd1755 : q <= 28'h0017d98; 
			12'd1756 : q <= 28'h0006485; 
			12'd1757 : q <= 28'h0008f7d; 
			12'd1758 : q <= 28'h000728e; 
			12'd1759 : q <= 28'h000628a; 
			12'd1760 : q <= 28'hfff9574; 
			12'd1761 : q <= 28'h0008b6c; 
			12'd1762 : q <= 28'hffc207e; 
			12'd1763 : q <= 28'h0027eb7; 
			12'd1764 : q <= 28'hfff6584; 
			12'd1765 : q <= 28'h0027d9b; 
			12'd1766 : q <= 28'hfff5381; 
			12'd1767 : q <= 28'hffc2885; 
			12'd1768 : q <= 28'h00477a9; 
			12'd1769 : q <= 28'h0018559; 
			12'd1770 : q <= 28'h0009373; 
			12'd1771 : q <= 28'h0007388; 
			12'd1772 : q <= 28'h0008b6e; 
			12'd1773 : q <= 28'h0008968; 
			12'd1774 : q <= 28'h0007290; 
			12'd1775 : q <= 28'hfff7387; 
			12'd1776 : q <= 28'h0008d70; 
			12'd1777 : q <= 28'h001843f; 
			12'd1778 : q <= 28'h0006283; 
			12'd1779 : q <= 28'h0007d98; 
			12'd1780 : q <= 28'h000bd7a; 
			12'd1781 : q <= 28'hffd5d86; 
			12'd1782 : q <= 28'h002825c; 
			12'd1783 : q <= 28'h003856e; 
			12'd1784 : q <= 28'h00176a2; 
			12'd1785 : q <= 28'h0009773; 
			12'd1786 : q <= 28'h0006386; 
			12'd1787 : q <= 28'h0008d74; 
			12'd1788 : q <= 28'h0007492; 
			12'd1789 : q <= 28'h0008875; 
			12'd1790 : q <= 28'h0006585; 
			12'd1791 : q <= 28'hffb4886; 
			12'd1792 : q <= 28'h0007597; 
			12'd1793 : q <= 28'h0058549; 
			12'd1794 : q <= 28'h000708c; 
			12'd1795 : q <= 28'hffa5084; 
			12'd1796 : q <= 28'hffd5281; 
			12'd1797 : q <= 28'hfffa37c; 
			12'd1798 : q <= 28'hffe4680; 
			12'd1799 : q <= 28'h0007795; 
			12'd1800 : q <= 28'h0008463; 
			12'd1801 : q <= 28'hffe3485; 
			12'd1802 : q <= 28'hffe9d76; 
			12'd1803 : q <= 28'h0018b70; 
			12'd1804 : q <= 28'h000a277; 
			12'd1805 : q <= 28'h0018766; 
			12'd1806 : q <= 28'h000708b; 
			12'd1807 : q <= 28'h000977c; 
			12'd1808 : q <= 28'h0006886; 
			12'd1809 : q <= 28'h006845e; 
			12'd1810 : q <= 28'hff4217f; 
			12'd1811 : q <= 28'h000a47c; 
			12'd1812 : q <= 28'hfe80c7e; 
			12'd1813 : q <= 28'h0007689; 
			12'd1814 : q <= 28'h000a076; 
			12'd1815 : q <= 28'h0008976; 
			12'd1816 : q <= 28'h0006183; 
			12'd1817 : q <= 28'h0007491; 
			12'd1818 : q <= 28'hffca878; 
			12'd1819 : q <= 28'h003854d; 
			12'd1820 : q <= 28'h0008569; 
			12'd1821 : q <= 28'hfffa27e; 
			12'd1822 : q <= 28'h0006183; 
			12'd1823 : q <= 28'h0017e9f; 
			12'd1824 : q <= 28'h0147e21; 
			12'd1825 : q <= 28'hfe7c180; 
			12'd1826 : q <= 28'h0005e83; 
			12'd1827 : q <= 28'hffcab7d; 
			12'd1828 : q <= 28'h0047f2f; 
			12'd1829 : q <= 28'h000758d; 
			12'd1830 : q <= 28'h0008362; 
			12'd1831 : q <= 28'hfff6f8b; 
			12'd1832 : q <= 28'h00d77af; 
			12'd1833 : q <= 28'h0006e87; 
			12'd1834 : q <= 28'h0008970; 
			12'd1835 : q <= 28'h01a8311; 
			12'd1836 : q <= 28'h0006986; 
			12'd1837 : q <= 28'h00c8a71; 
			12'd1838 : q <= 28'h0006f8a; 
			12'd1839 : q <= 28'hffa9980; 
			12'd1840 : q <= 28'h00d7e23; 
			12'd1841 : q <= 28'hffda37f; 
			12'd1842 : q <= 28'hfdb197e; 
			12'd1843 : q <= 28'hffc5485; 
			12'd1844 : q <= 28'h000708a; 
			12'd1845 : q <= 28'hfff4784; 
			12'd1846 : q <= 28'hfffb279; 
			12'd1847 : q <= 28'h0007fa1; 
			12'd1848 : q <= 28'hfff4c80; 
			12'd1849 : q <= 28'h0008762; 
			12'd1850 : q <= 28'hffe347f; 
			12'd1851 : q <= 28'h00780b1; 
			12'd1852 : q <= 28'h02b7e25; 
			12'd1853 : q <= 28'h0008f7b; 
			12'd1854 : q <= 28'h0008569; 
			12'd1855 : q <= 28'h05c8560; 
			12'd1856 : q <= 28'hffe9a76; 
			12'd1857 : q <= 28'hfff6888; 
			12'd1858 : q <= 28'h0007597; 
			12'd1859 : q <= 28'h0008a6f; 
			12'd1860 : q <= 28'h0008567; 
			12'd1861 : q <= 28'h000768e; 
			12'd1862 : q <= 28'hfff9e77; 
			12'd1863 : q <= 28'hfffaf80; 
			12'd1864 : q <= 28'h0006f89; 
			12'd1865 : q <= 28'h0007992; 
			12'd1866 : q <= 28'h002825d; 
			12'd1867 : q <= 28'h0008e75; 
			12'd1868 : q <= 28'h000896f; 
			12'd1869 : q <= 28'h000718b; 
			12'd1870 : q <= 28'h0006784; 
			12'd1871 : q <= 28'h0017e90; 
			12'd1872 : q <= 28'hffbcc7a; 
			12'd1873 : q <= 28'hffd6584; 
			12'd1874 : q <= 28'hff6057e; 
			12'd1875 : q <= 28'h0006688; 
			12'd1876 : q <= 28'h0017696; 
			12'd1877 : q <= 28'hfffa680; 
			12'd1878 : q <= 28'h0188669; 
			12'd1879 : q <= 28'h0017c96; 
			12'd1880 : q <= 28'h0006484; 
			12'd1881 : q <= 28'h000957f; 
			12'd1882 : q <= 28'hffa207e; 
			12'd1883 : q <= 28'hfff9280; 
			12'd1884 : q <= 28'h001866c; 
			12'd1885 : q <= 28'h0007194; 
			12'd1886 : q <= 28'h0009373; 
			12'd1887 : q <= 28'hffd3084; 
			12'd1888 : q <= 28'hfffa879; 
			12'd1889 : q <= 28'h0018655; 
			12'd1890 : q <= 28'h000896d; 
			12'd1891 : q <= 28'h0018094; 
			12'd1892 : q <= 28'h00179aa; 
			12'd1893 : q <= 28'h000896e; 
			12'd1894 : q <= 28'h0057f30; 
			12'd1895 : q <= 28'h0017e94; 
			12'd1896 : q <= 28'h0028569; 
			12'd1897 : q <= 28'h0008c7a; 
			12'd1898 : q <= 28'h000789a; 
			12'd1899 : q <= 28'h001844e; 
			12'd1900 : q <= 28'h000856a; 
			12'd1901 : q <= 28'h000967b; 
			12'd1902 : q <= 28'hffe2c7f; 
			12'd1903 : q <= 28'h0006f85; 
			12'd1904 : q <= 28'h00079b0; 
			12'd1905 : q <= 28'h000866f; 
			12'd1906 : q <= 28'h0017ac8; 
			12'd1907 : q <= 28'h0006989; 
			12'd1908 : q <= 28'h00179a4; 
			12'd1909 : q <= 28'hffe3f84; 
			12'd1910 : q <= 28'hffc9376; 
			12'd1911 : q <= 28'h0018452; 
			12'd1912 : q <= 28'hfff6383; 
			12'd1913 : q <= 28'h0017ca1; 
			12'd1914 : q <= 28'h000835f; 
			12'd1915 : q <= 28'hffb917d; 
			12'd1916 : q <= 28'h0004180; 
			12'd1917 : q <= 28'h0017b91; 
			12'd1918 : q <= 28'h0067f2d; 
			12'd1919 : q <= 28'h0007e8c; 
			12'd1920 : q <= 28'h0088047; 
			12'd1921 : q <= 28'hffdb47f; 
			12'd1922 : q <= 28'h0008360; 
			12'd1923 : q <= 28'hfe8a566; 
			12'd1924 : q <= 28'h0016693; 
			12'd1925 : q <= 28'h0005b8d; 
			12'd1926 : q <= 28'h0006c89; 
			12'd1927 : q <= 28'h0005e8f; 
			12'd1928 : q <= 28'h0008b66; 
			12'd1929 : q <= 28'h0008654; 
			12'd1930 : q <= 28'hffe6e87; 
			12'd1931 : q <= 28'h00273a5; 
			12'd1932 : q <= 28'h0006e89; 
			12'd1933 : q <= 28'h0008861; 
			12'd1934 : q <= 28'h0006e89; 
			12'd1935 : q <= 28'h0006c8d; 
			12'd1936 : q <= 28'h0128744; 
			12'd1937 : q <= 28'h0005b85; 
			12'd1938 : q <= 28'h0108549; 
			12'd1939 : q <= 28'h0005c85; 
			12'd1940 : q <= 28'h0008c65; 
			12'd1941 : q <= 28'h0005f85; 
			12'd1942 : q <= 28'h0009675; 
			12'd1943 : q <= 28'h0006889; 
			12'd1944 : q <= 28'h0006087; 
			12'd1945 : q <= 28'hfe74b81; 
			12'd1946 : q <= 28'h0007cac; 
			12'd1947 : q <= 28'h0006f8e; 
			12'd1948 : q <= 28'hff85087; 
			12'd1949 : q <= 28'hfffa776; 
			12'd1950 : q <= 28'h0048450; 
			12'd1951 : q <= 28'h0006888; 
			12'd1952 : q <= 28'h0017fa9; 
			12'd1953 : q <= 28'h0009773; 
			12'd1954 : q <= 28'h000885c; 
			12'd1955 : q <= 28'hfff3b7f; 
			12'd1956 : q <= 28'h0009677; 
			12'd1957 : q <= 28'h0027f30; 
			12'd1958 : q <= 28'h000967a; 
			12'd1959 : q <= 28'h0008359; 
			12'd1960 : q <= 28'h0008869; 
			12'd1961 : q <= 28'h0006e8a; 
			12'd1962 : q <= 28'hff84484; 
			12'd1963 : q <= 28'h0047f3b; 
			12'd1964 : q <= 28'h0008d76; 
			12'd1965 : q <= 28'h0009072; 
			12'd1966 : q <= 28'hffeab7e; 
			12'd1967 : q <= 28'h0008664; 
			12'd1968 : q <= 28'h0007a8c; 
			12'd1969 : q <= 28'hfffb178; 
			12'd1970 : q <= 28'hfff688c; 
			12'd1971 : q <= 28'hfff5481; 
			12'd1972 : q <= 28'h0007fa3; 
			12'd1973 : q <= 28'h001779f; 
			12'd1974 : q <= 28'hffa3b85; 
			12'd1975 : q <= 28'hffb1e7e; 
			12'd1976 : q <= 28'h0008869; 
			12'd1977 : q <= 28'hffca077; 
			12'd1978 : q <= 28'hffe5786; 
			12'd1979 : q <= 28'h0005c82; 
			12'd1980 : q <= 28'h0017d9e; 
			12'd1981 : q <= 28'hfff4380; 
			12'd1982 : q <= 28'h0006f90; 
			12'd1983 : q <= 28'hff5a678; 
			12'd1984 : q <= 28'hffb6187; 
			12'd1985 : q <= 28'hffb5281; 
			12'd1986 : q <= 28'h0018472; 
			12'd1987 : q <= 28'h0006686; 
			12'd1988 : q <= 28'h000a17d; 
			12'd1989 : q <= 28'h00078a6; 
			12'd1990 : q <= 28'hfff5d85; 
			12'd1991 : q <= 28'h0008463; 
			12'd1992 : q <= 28'hfffbc80; 
			12'd1993 : q <= 28'h000718c; 
			12'd1994 : q <= 28'h000987c; 
			12'd1995 : q <= 28'h0009870; 
			12'd1996 : q <= 28'h0008875; 
			12'd1997 : q <= 28'h001814b; 
			12'd1998 : q <= 28'hffa4185; 
			12'd1999 : q <= 28'h000718c; 
			12'd2000 : q <= 28'h0008868; 
			12'd2001 : q <= 28'h0006886; 
			12'd2002 : q <= 28'h000917d; 
			12'd2003 : q <= 28'h0006986; 
			12'd2004 : q <= 28'h00181bb; 
			12'd2005 : q <= 28'h0009975; 
			12'd2006 : q <= 28'hffa6a87; 
			12'd2007 : q <= 28'h0008f73; 
			12'd2008 : q <= 28'h0006889; 
			12'd2009 : q <= 28'h0006f8b; 
			12'd2010 : q <= 28'hffd2a83; 
			12'd2011 : q <= 28'h0027f30; 
			12'd2012 : q <= 28'h0007c9c; 
			12'd2013 : q <= 28'hfffa078; 
			12'd2014 : q <= 28'h0008e67; 
			12'd2015 : q <= 28'h0006986; 
			12'd2016 : q <= 28'h0017991; 
			12'd2017 : q <= 28'h0077f2c; 
			12'd2018 : q <= 28'h000896f; 
			12'd2019 : q <= 28'h000896f; 
			12'd2020 : q <= 28'hfff5784; 
			12'd2021 : q <= 28'h00b7aba; 
			12'd2022 : q <= 28'h0008090; 
			12'd2023 : q <= 28'h0006684; 
			12'd2024 : q <= 28'h000688a; 
			12'd2025 : q <= 28'hfff6886; 
			12'd2026 : q <= 28'h0007da3; 
			12'd2027 : q <= 28'h001804b; 
			12'd2028 : q <= 28'h0027ea1; 
			12'd2029 : q <= 28'h000886d; 
			12'd2030 : q <= 28'h0007f98; 
			12'd2031 : q <= 28'h0007595; 
			12'd2032 : q <= 28'h0007595; 
			12'd2033 : q <= 28'h0006585; 
			12'd2034 : q <= 28'h000947d; 
			12'd2035 : q <= 28'h0006f8c; 
			12'd2036 : q <= 28'h0008962; 
			12'd2037 : q <= 28'h0018048; 
			12'd2038 : q <= 28'hfed1f83; 
			12'd2039 : q <= 28'h00679b3; 
			12'd2040 : q <= 28'h0008b77; 
			12'd2041 : q <= 28'h0006784; 
			12'd2042 : q <= 28'h0006e84; 
			12'd2043 : q <= 28'h0009f78; 
			12'd2044 : q <= 28'h0008971; 
			12'd2045 : q <= 28'h000876c; 
			12'd2046 : q <= 28'hffd4284; 
			12'd2047 : q <= 28'h0057ac2; 
			12'd2048 : q <= 28'h0008877; 
			12'd2049 : q <= 28'h0037f25; 
			12'd2050 : q <= 28'hff4a480; 
			12'd2051 : q <= 28'h0047391; 
			12'd2052 : q <= 28'hffc4683; 
			12'd2053 : q <= 28'h0008361; 
			12'd2054 : q <= 28'h01081a8; 
			12'd2055 : q <= 28'h0008566; 
			12'd2056 : q <= 28'h0007f98; 
			12'd2057 : q <= 28'hffc6084; 
			12'd2058 : q <= 28'h000a981; 
			12'd2059 : q <= 28'h0137ace; 
			12'd2060 : q <= 28'h0017e92; 
			12'd2061 : q <= 28'hfee0d7e; 
			12'd2062 : q <= 28'h08a831d; 
			12'd2063 : q <= 28'h0007391; 
			12'd2064 : q <= 28'h000896b; 
			12'd2065 : q <= 28'h0009776; 
			12'd2066 : q <= 28'h0008670; 
			12'd2067 : q <= 28'h0006784; 
			12'd2068 : q <= 28'hffabe82; 
			12'd2069 : q <= 28'h0005481; 
			12'd2070 : q <= 28'h0017c94; 
			12'd2071 : q <= 28'hff56e89; 
			12'd2072 : q <= 28'h027852b; 
			12'd2073 : q <= 28'h00379ac; 
			12'd2074 : q <= 28'h000957a; 
			12'd2075 : q <= 28'h0017f3b; 
			12'd2076 : q <= 28'hffd7986; 
			12'd2077 : q <= 28'h001815b; 
			12'd2078 : q <= 28'h0007c8f; 
			12'd2079 : q <= 28'h00279ad; 
			12'd2080 : q <= 28'h000876d; 
			12'd2081 : q <= 28'h000738d; 
			12'd2082 : q <= 28'hfff6a8b; 
			12'd2083 : q <= 28'h00178a6; 
			12'd2084 : q <= 28'hffd3784; 
			12'd2085 : q <= 28'h000886e; 
			12'd2086 : q <= 28'h000758e; 
			12'd2087 : q <= 28'h0047e12; 
			12'd2088 : q <= 28'hff8b37f; 
			12'd2089 : q <= 28'h000728c; 
			12'd2090 : q <= 28'h0007888; 
			12'd2091 : q <= 28'h0006e88; 
			12'd2092 : q <= 28'hffb4385; 
			12'd2093 : q <= 28'h000856a; 
			12'd2094 : q <= 28'hff9a280; 
			12'd2095 : q <= 28'h0018159; 
			12'd2096 : q <= 28'h0057fb2; 
			12'd2097 : q <= 28'hffe5481; 
			12'd2098 : q <= 28'h0047fbb; 
			12'd2099 : q <= 28'h0006484; 
			12'd2100 : q <= 28'h000907e; 
			12'd2101 : q <= 28'h0009574; 
			12'd2102 : q <= 28'h0006d8b; 
			12'd2103 : q <= 28'h0008363; 
			12'd2104 : q <= 28'hffe9a7f; 
			12'd2105 : q <= 28'hffd4280; 
			12'd2106 : q <= 28'h0007c8e; 
			12'd2107 : q <= 28'h0009776; 
			12'd2108 : q <= 28'hffc5084; 
			12'd2109 : q <= 28'h0018158; 
			12'd2110 : q <= 28'h0007a96; 
			12'd2111 : q <= 28'h0006e89; 
			12'd2112 : q <= 28'h0008b76; 
			12'd2113 : q <= 28'h00279ad; 
			12'd2114 : q <= 28'h0006c8a; 
			12'd2115 : q <= 28'hfff9c77; 
			12'd2116 : q <= 28'h0009171; 
			12'd2117 : q <= 28'h0006084; 
			12'd2118 : q <= 28'h0007893; 
			12'd2119 : q <= 28'h000728f; 
			12'd2120 : q <= 28'h0008b64; 
			12'd2121 : q <= 28'h0007490; 
			12'd2122 : q <= 28'h0009378; 
			12'd2123 : q <= 28'h0008460; 
			12'd2124 : q <= 28'h001809d; 
			12'd2125 : q <= 28'h0008a70; 
			12'd2126 : q <= 28'h00b8434; 
			12'd2127 : q <= 28'h0006383; 
			12'd2128 : q <= 28'h0007d8a; 
			12'd2129 : q <= 28'hffcb27a; 
			12'd2130 : q <= 28'h035854d; 
			12'd2131 : q <= 28'h0008a72; 
			12'd2132 : q <= 28'h0007b9a; 
			12'd2133 : q <= 28'hfff6584; 
			12'd2134 : q <= 28'h0028b6b; 
			12'd2135 : q <= 28'h00b79a6;
			default	 : q <= 28'h0000000;
		endcase	
	end
	assign out = q;
endmodule