
module classifier_tb;

    reg clk;
    reg rst;
    reg en;
    reg[20*20*9 - 1 : 0] image;
    wire face_status;
    wire request_new_data;

    top_level_classifier#(.WIDTH(20), .BITSIZE(9))
    toplevel (
        .clk(clk),
        .rst(rst),
        .en(en),
        .image(image),
        .face_status(face_status),
        .request_new_data(request_new_data)
    );

    initial begin
        clk = 1'b0;
        rst = 1'b1;
        en = 1'b0;

        image[8 : 0] = 9'd0;
        image[17 : 9] = 9'd1;
        image[26 : 18] = 9'd1;
        image[35 : 27] = 9'd1;
        image[44 : 36] = 9'd2;
        image[53 : 45] = 9'd3;
        image[62 : 54] = 9'd4;
        image[71 : 63] = 9'd5;
        image[80 : 72] = 9'd6;
        image[89 : 81] = 9'd7;
        image[98 : 90] = 9'd8;
        image[107 : 99] = 9'd9;
        image[116 : 108] = 9'd10;
        image[125 : 117] = 9'd11;
        image[134 : 126] = 9'd12;
        image[143 : 135] = 9'd13;
        image[152 : 144] = 9'd13;
        image[161 : 153] = 9'd14;
        image[170 : 162] = 9'd15;
        image[179 : 171] = 9'd16;
        image[188 : 180] = 9'd0;
        image[197 : 189] = 9'd2;
        image[206 : 198] = 9'd2;
        image[215 : 207] = 9'd2;
        image[224 : 216] = 9'd4;
        image[233 : 225] = 9'd6;
        image[242 : 234] = 9'd8;
        image[251 : 243] = 9'd10;
        image[260 : 252] = 9'd12;
        image[269 : 261] = 9'd14;
        image[278 : 270] = 9'd16;
        image[287 : 279] = 9'd18;
        image[296 : 288] = 9'd20;
        image[305 : 297] = 9'd22;
        image[314 : 306] = 9'd24;
        image[323 : 315] = 9'd25;
        image[332 : 324] = 9'd25;
        image[341 : 333] = 9'd27;
        image[350 : 342] = 9'd29;
        image[359 : 351] = 9'd31;
        image[368 : 360] = 9'd0;
        image[377 : 369] = 9'd2;
        image[386 : 378] = 9'd2;
        image[395 : 387] = 9'd2;
        image[404 : 396] = 9'd5;
        image[413 : 405] = 9'd8;
        image[422 : 414] = 9'd11;
        image[431 : 423] = 9'd14;
        image[440 : 432] = 9'd17;
        image[449 : 441] = 9'd20;
        image[458 : 450] = 9'd23;
        image[467 : 459] = 9'd26;
        image[476 : 468] = 9'd29;
        image[485 : 477] = 9'd32;
        image[494 : 486] = 9'd35;
        image[503 : 495] = 9'd37;
        image[512 : 504] = 9'd37;
        image[521 : 513] = 9'd40;
        image[530 : 522] = 9'd43;
        image[539 : 531] = 9'd46;
        image[548 : 540] = 9'd0;
        image[557 : 549] = 9'd2;
        image[566 : 558] = 9'd2;
        image[575 : 567] = 9'd2;
        image[584 : 576] = 9'd6;
        image[593 : 585] = 9'd10;
        image[602 : 594] = 9'd14;
        image[611 : 603] = 9'd18;
        image[620 : 612] = 9'd22;
        image[629 : 621] = 9'd26;
        image[638 : 630] = 9'd30;
        image[647 : 639] = 9'd34;
        image[656 : 648] = 9'd38;
        image[665 : 657] = 9'd42;
        image[674 : 666] = 9'd46;
        image[683 : 675] = 9'd49;
        image[692 : 684] = 9'd50;
        image[701 : 693] = 9'd53;
        image[710 : 702] = 9'd57;
        image[719 : 711] = 9'd61;
        image[728 : 720] = 9'd0;
        image[737 : 729] = 9'd2;
        image[746 : 738] = 9'd2;
        image[755 : 747] = 9'd3;
        image[764 : 756] = 9'd8;
        image[773 : 765] = 9'd13;
        image[782 : 774] = 9'd18;
        image[791 : 783] = 9'd23;
        image[800 : 792] = 9'd28;
        image[809 : 801] = 9'd33;
        image[818 : 810] = 9'd38;
        image[827 : 819] = 9'd43;
        image[836 : 828] = 9'd48;
        image[845 : 837] = 9'd53;
        image[854 : 846] = 9'd58;
        image[863 : 855] = 9'd62;
        image[872 : 864] = 9'd64;
        image[881 : 873] = 9'd67;
        image[890 : 882] = 9'd71;
        image[899 : 891] = 9'd76;
        image[908 : 900] = 9'd0;
        image[917 : 909] = 9'd2;
        image[926 : 918] = 9'd2;
        image[935 : 927] = 9'd3;
        image[944 : 936] = 9'd9;
        image[953 : 945] = 9'd15;
        image[962 : 954] = 9'd21;
        image[971 : 963] = 9'd27;
        image[980 : 972] = 9'd33;
        image[989 : 981] = 9'd39;
        image[998 : 990] = 9'd45;
        image[1007 : 999] = 9'd51;
        image[1016 : 1008] = 9'd57;
        image[1025 : 1017] = 9'd63;
        image[1034 : 1026] = 9'd69;
        image[1043 : 1035] = 9'd74;
        image[1052 : 1044] = 9'd77;
        image[1061 : 1053] = 9'd80;
        image[1070 : 1062] = 9'd84;
        image[1079 : 1071] = 9'd89;
        image[1088 : 1080] = 9'd0;
        image[1097 : 1089] = 9'd2;
        image[1106 : 1098] = 9'd2;
        image[1115 : 1107] = 9'd3;
        image[1124 : 1116] = 9'd10;
        image[1133 : 1125] = 9'd16;
        image[1142 : 1134] = 9'd22;
        image[1151 : 1143] = 9'd29;
        image[1160 : 1152] = 9'd36;
        image[1169 : 1161] = 9'd43;
        image[1178 : 1170] = 9'd50;
        image[1187 : 1179] = 9'd57;
        image[1196 : 1188] = 9'd64;
        image[1205 : 1197] = 9'd70;
        image[1214 : 1206] = 9'd76;
        image[1223 : 1215] = 9'd82;
        image[1232 : 1224] = 9'd86;
        image[1241 : 1233] = 9'd89;
        image[1250 : 1242] = 9'd93;
        image[1259 : 1251] = 9'd98;
        image[1268 : 1260] = 9'd0;
        image[1277 : 1269] = 9'd2;
        image[1286 : 1278] = 9'd2;
        image[1295 : 1287] = 9'd3;
        image[1304 : 1296] = 9'd10;
        image[1313 : 1305] = 9'd16;
        image[1322 : 1314] = 9'd22;
        image[1331 : 1323] = 9'd29;
        image[1340 : 1332] = 9'd36;
        image[1349 : 1341] = 9'd44;
        image[1358 : 1350] = 9'd52;
        image[1367 : 1359] = 9'd60;
        image[1376 : 1368] = 9'd67;
        image[1385 : 1377] = 9'd73;
        image[1394 : 1386] = 9'd79;
        image[1403 : 1395] = 9'd85;
        image[1412 : 1404] = 9'd90;
        image[1421 : 1413] = 9'd93;
        image[1430 : 1422] = 9'd97;
        image[1439 : 1431] = 9'd102;
        image[1448 : 1440] = 9'd0;
        image[1457 : 1449] = 9'd2;
        image[1466 : 1458] = 9'd2;
        image[1475 : 1467] = 9'd3;
        image[1484 : 1476] = 9'd10;
        image[1493 : 1485] = 9'd16;
        image[1502 : 1494] = 9'd22;
        image[1511 : 1503] = 9'd30;
        image[1520 : 1512] = 9'd37;
        image[1529 : 1521] = 9'd46;
        image[1538 : 1530] = 9'd55;
        image[1547 : 1539] = 9'd64;
        image[1556 : 1548] = 9'd72;
        image[1565 : 1557] = 9'd79;
        image[1574 : 1566] = 9'd86;
        image[1583 : 1575] = 9'd93;
        image[1592 : 1584] = 9'd99;
        image[1601 : 1593] = 9'd103;
        image[1610 : 1602] = 9'd107;
        image[1619 : 1611] = 9'd112;
        image[1628 : 1620] = 9'd0;
        image[1637 : 1629] = 9'd2;
        image[1646 : 1638] = 9'd2;
        image[1655 : 1647] = 9'd3;
        image[1664 : 1656] = 9'd11;
        image[1673 : 1665] = 9'd18;
        image[1682 : 1674] = 9'd25;
        image[1691 : 1683] = 9'd34;
        image[1700 : 1692] = 9'd41;
        image[1709 : 1701] = 9'd51;
        image[1718 : 1710] = 9'd61;
        image[1727 : 1719] = 9'd71;
        image[1736 : 1728] = 9'd80;
        image[1745 : 1737] = 9'd88;
        image[1754 : 1746] = 9'd96;
        image[1763 : 1755] = 9'd104;
        image[1772 : 1764] = 9'd111;
        image[1781 : 1773] = 9'd116;
        image[1790 : 1782] = 9'd120;
        image[1799 : 1791] = 9'd125;
        image[1808 : 1800] = 9'd0;
        image[1817 : 1809] = 9'd2;
        image[1826 : 1818] = 9'd2;
        image[1835 : 1827] = 9'd3;
        image[1844 : 1836] = 9'd12;
        image[1853 : 1845] = 9'd20;
        image[1862 : 1854] = 9'd28;
        image[1871 : 1863] = 9'd38;
        image[1880 : 1872] = 9'd45;
        image[1889 : 1881] = 9'd56;
        image[1898 : 1890] = 9'd67;
        image[1907 : 1899] = 9'd78;
        image[1916 : 1908] = 9'd88;
        image[1925 : 1917] = 9'd97;
        image[1934 : 1926] = 9'd106;
        image[1943 : 1935] = 9'd115;
        image[1952 : 1944] = 9'd123;
        image[1961 : 1953] = 9'd129;
        image[1970 : 1962] = 9'd133;
        image[1979 : 1971] = 9'd138;
        image[1988 : 1980] = 9'd0;
        image[1997 : 1989] = 9'd2;
        image[2006 : 1998] = 9'd2;
        image[2015 : 2007] = 9'd3;
        image[2024 : 2016] = 9'd13;
        image[2033 : 2025] = 9'd22;
        image[2042 : 2034] = 9'd31;
        image[2051 : 2043] = 9'd42;
        image[2060 : 2052] = 9'd49;
        image[2069 : 2061] = 9'd61;
        image[2078 : 2070] = 9'd73;
        image[2087 : 2079] = 9'd85;
        image[2096 : 2088] = 9'd96;
        image[2105 : 2097] = 9'd106;
        image[2114 : 2106] = 9'd116;
        image[2123 : 2115] = 9'd126;
        image[2132 : 2124] = 9'd135;
        image[2141 : 2133] = 9'd142;
        image[2150 : 2142] = 9'd146;
        image[2159 : 2151] = 9'd151;
        image[2168 : 2160] = 9'd0;
        image[2177 : 2169] = 9'd2;
        image[2186 : 2178] = 9'd2;
        image[2195 : 2187] = 9'd3;
        image[2204 : 2196] = 9'd14;
        image[2213 : 2205] = 9'd24;
        image[2222 : 2214] = 9'd34;
        image[2231 : 2223] = 9'd45;
        image[2240 : 2232] = 9'd52;
        image[2249 : 2241] = 9'd65;
        image[2258 : 2250] = 9'd78;
        image[2267 : 2259] = 9'd91;
        image[2276 : 2268] = 9'd103;
        image[2285 : 2277] = 9'd114;
        image[2294 : 2286] = 9'd125;
        image[2303 : 2295] = 9'd136;
        image[2312 : 2304] = 9'd146;
        image[2321 : 2313] = 9'd153;
        image[2330 : 2322] = 9'd157;
        image[2339 : 2331] = 9'd162;
        image[2348 : 2340] = 9'd0;
        image[2357 : 2349] = 9'd2;
        image[2366 : 2358] = 9'd2;
        image[2375 : 2367] = 9'd3;
        image[2384 : 2376] = 9'd14;
        image[2393 : 2385] = 9'd25;
        image[2402 : 2394] = 9'd36;
        image[2411 : 2403] = 9'd47;
        image[2420 : 2412] = 9'd54;
        image[2429 : 2421] = 9'd68;
        image[2438 : 2430] = 9'd82;
        image[2447 : 2439] = 9'd96;
        image[2456 : 2448] = 9'd109;
        image[2465 : 2457] = 9'd121;
        image[2474 : 2466] = 9'd133;
        image[2483 : 2475] = 9'd145;
        image[2492 : 2484] = 9'd156;
        image[2501 : 2493] = 9'd163;
        image[2510 : 2502] = 9'd167;
        image[2519 : 2511] = 9'd172;
        image[2528 : 2520] = 9'd0;
        image[2537 : 2529] = 9'd2;
        image[2546 : 2538] = 9'd2;
        image[2555 : 2547] = 9'd3;
        image[2564 : 2556] = 9'd14;
        image[2573 : 2565] = 9'd26;
        image[2582 : 2574] = 9'd38;
        image[2591 : 2583] = 9'd49;
        image[2600 : 2592] = 9'd56;
        image[2609 : 2601] = 9'd71;
        image[2618 : 2610] = 9'd86;
        image[2627 : 2619] = 9'd101;
        image[2636 : 2628] = 9'd115;
        image[2645 : 2637] = 9'd128;
        image[2654 : 2646] = 9'd141;
        image[2663 : 2655] = 9'd154;
        image[2672 : 2664] = 9'd166;
        image[2681 : 2673] = 9'd173;
        image[2690 : 2682] = 9'd177;
        image[2699 : 2691] = 9'd182;
        image[2708 : 2700] = 9'd0;
        image[2717 : 2709] = 9'd2;
        image[2726 : 2718] = 9'd2;
        image[2735 : 2727] = 9'd3;
        image[2744 : 2736] = 9'd14;
        image[2753 : 2745] = 9'd27;
        image[2762 : 2754] = 9'd40;
        image[2771 : 2763] = 9'd51;
        image[2780 : 2772] = 9'd58;
        image[2789 : 2781] = 9'd74;
        image[2798 : 2790] = 9'd90;
        image[2807 : 2799] = 9'd106;
        image[2816 : 2808] = 9'd121;
        image[2825 : 2817] = 9'd135;
        image[2834 : 2826] = 9'd149;
        image[2843 : 2835] = 9'd163;
        image[2852 : 2844] = 9'd175;
        image[2861 : 2853] = 9'd182;
        image[2870 : 2862] = 9'd186;
        image[2879 : 2871] = 9'd191;
        image[2888 : 2880] = 9'd0;
        image[2897 : 2889] = 9'd2;
        image[2906 : 2898] = 9'd2;
        image[2915 : 2907] = 9'd3;
        image[2924 : 2916] = 9'd14;
        image[2933 : 2925] = 9'd27;
        image[2942 : 2934] = 9'd41;
        image[2951 : 2943] = 9'd53;
        image[2960 : 2952] = 9'd60;
        image[2969 : 2961] = 9'd76;
        image[2978 : 2970] = 9'd93;
        image[2987 : 2979] = 9'd110;
        image[2996 : 2988] = 9'd126;
        image[3005 : 2997] = 9'd141;
        image[3014 : 3006] = 9'd156;
        image[3023 : 3015] = 9'd171;
        image[3032 : 3024] = 9'd183;
        image[3041 : 3033] = 9'd190;
        image[3050 : 3042] = 9'd194;
        image[3059 : 3051] = 9'd199;
        image[3068 : 3060] = 9'd0;
        image[3077 : 3069] = 9'd2;
        image[3086 : 3078] = 9'd2;
        image[3095 : 3087] = 9'd3;
        image[3104 : 3096] = 9'd14;
        image[3113 : 3105] = 9'd27;
        image[3122 : 3114] = 9'd41;
        image[3131 : 3123] = 9'd54;
        image[3140 : 3132] = 9'd62;
        image[3149 : 3141] = 9'd79;
        image[3158 : 3150] = 9'd97;
        image[3167 : 3159] = 9'd115;
        image[3176 : 3168] = 9'd132;
        image[3185 : 3177] = 9'd148;
        image[3194 : 3186] = 9'd164;
        image[3203 : 3195] = 9'd179;
        image[3212 : 3204] = 9'd191;
        image[3221 : 3213] = 9'd198;
        image[3230 : 3222] = 9'd202;
        image[3239 : 3231] = 9'd207;
        image[3248 : 3240] = 9'd0;
        image[3257 : 3249] = 9'd2;
        image[3266 : 3258] = 9'd2;
        image[3275 : 3267] = 9'd3;
        image[3284 : 3276] = 9'd14;
        image[3293 : 3285] = 9'd27;
        image[3302 : 3294] = 9'd41;
        image[3311 : 3303] = 9'd54;
        image[3320 : 3312] = 9'd63;
        image[3329 : 3321] = 9'd81;
        image[3338 : 3330] = 9'd100;
        image[3347 : 3339] = 9'd119;
        image[3356 : 3348] = 9'd137;
        image[3365 : 3357] = 9'd154;
        image[3374 : 3366] = 9'd171;
        image[3383 : 3375] = 9'd186;
        image[3392 : 3384] = 9'd198;
        image[3401 : 3393] = 9'd205;
        image[3410 : 3402] = 9'd209;
        image[3419 : 3411] = 9'd214;
        image[3428 : 3420] = 9'd0;
        image[3437 : 3429] = 9'd2;
        image[3446 : 3438] = 9'd2;
        image[3455 : 3447] = 9'd3;
        image[3464 : 3456] = 9'd14;
        image[3473 : 3465] = 9'd27;
        image[3482 : 3474] = 9'd41;
        image[3491 : 3483] = 9'd54;
        image[3500 : 3492] = 9'd64;
        image[3509 : 3501] = 9'd83;
        image[3518 : 3510] = 9'd103;
        image[3527 : 3519] = 9'd123;
        image[3536 : 3528] = 9'd142;
        image[3545 : 3537] = 9'd160;
        image[3554 : 3546] = 9'd177;
        image[3563 : 3555] = 9'd192;
        image[3572 : 3564] = 9'd204;
        image[3581 : 3573] = 9'd211;
        image[3590 : 3582] = 9'd215;
        image[3599 : 3591] = 9'd220;

        #15
        rst = 1'b0;
        en = 1'b1;  
    end

    always #5 clk = !clk;
endmodule 