module rect2_rom(
	input [11:0] addr,
	input clk,
	output[22:0] out
);
	reg[22:0] q;

	always @(posedge clk)
	begin
		case(addr)
			12'd1    : q <= 23'h21a5c2;
			12'd2    : q <= 23'h3388c4;
			12'd3    : q <= 23'h30a9e3;
			12'd4    : q <= 23'h22a443;
			12'd5    : q <= 23'h349443;
			12'd6    : q <= 23'h320d83;
			12'd7    : q <= 23'h233544;
			12'd8    : q <= 23'h21a9c4;
			12'd9    : q <= 23'h27046a;
			12'd10   : q <= 23'h33b0a4;
			12'd11   : q <= 23'h3384c3;
			12'd12   : q <= 23'h20a621;
			12'd13   : q <= 23'h281c81;
			12'd14   : q <= 23'h22c841;
			12'd15   : q <= 23'h27086c;
			12'd16   : q <= 23'h220046;
			12'd17   : q <= 23'h342cc8;
			12'd18   : q <= 23'h22a141;
			12'd19   : q <= 23'h37b0a1;
			12'd20   : q <= 23'h329943;
			12'd21   : q <= 23'h24ac47;
			12'd22   : q <= 23'h31a484;
			12'd23   : q <= 23'h341485;
			12'd24   : q <= 23'h22a944;
			12'd25   : q <= 23'h340cc3;
			12'd26   : q <= 23'h24c024;
			12'd27   : q <= 23'h302682;
			12'd28   : q <= 23'h348051;
			12'd29   : q <= 23'h358044;
			12'd30   : q <= 23'h338444;
			12'd31   : q <= 23'h370450;
			12'd32   : q <= 23'h201524;
			12'd33   : q <= 23'h26bca2;
			12'd34   : q <= 23'h218444;
			12'd35   : q <= 23'h2518e5;
			12'd36   : q <= 23'h320450;
			12'd37   : q <= 23'h204e81;
			12'd38   : q <= 23'h343881;
			12'd39   : q <= 23'h34bc41;
			12'd40   : q <= 23'h303922;
			12'd41   : q <= 23'h22a462;
			12'd42   : q <= 23'h24ac48;
			12'd43   : q <= 23'h21a9a4;
			12'd44   : q <= 23'h260c82;
			12'd45   : q <= 23'h343084;
			12'd46   : q <= 23'h278c83;
			12'd47   : q <= 23'h348453;
			12'd48   : q <= 23'h358044;
			12'd49   : q <= 23'h330463;
			12'd50   : q <= 23'h26bca2;
			12'd51   : q <= 23'h218c6a;
			12'd52   : q <= 23'h31a5e5;
			12'd53   : q <= 23'h331d02;
			12'd54   : q <= 23'h2510c5;
			12'd55   : q <= 23'h241044;
			12'd56   : q <= 23'h27b021;
			12'd57   : q <= 23'h21b041;
			12'd58   : q <= 23'h383021;
			12'd59   : q <= 23'h21bc62;
			12'd60   : q <= 23'h232101;
			12'd61   : q <= 23'h31b021;
			12'd62   : q <= 23'h230581;
			12'd63   : q <= 23'h34bc41;
			12'd64   : q <= 23'h23c0c1;
			12'd65   : q <= 23'h301c82;
			12'd66   : q <= 23'h343082;
			12'd67   : q <= 23'h331823;
			12'd68   : q <= 23'h35c422;
			12'd69   : q <= 23'h24a841;
			12'd70   : q <= 23'h349844;
			12'd71   : q <= 23'h344422;
			12'd72   : q <= 23'h35c423;
			12'd73   : q <= 23'h243461;
			12'd74   : q <= 23'h358c42;
			12'd75   : q <= 23'h21b5c2;
			12'd76   : q <= 23'h252922;
			12'd77   : q <= 23'h302c61;
			12'd78   : q <= 23'h358446;
			12'd79   : q <= 23'h349c26;
			12'd80   : q <= 23'h308e43;
			12'd81   : q <= 23'h263443;
			12'd82   : q <= 23'h202664;
			12'd83   : q <= 23'h348049;
			12'd84   : q <= 23'h338c41;
			12'd85   : q <= 23'h368c41;
			12'd86   : q <= 23'h22b483;
			12'd87   : q <= 23'h368c41;
			12'd88   : q <= 23'h321982;
			12'd89   : q <= 23'h37b842;
			12'd90   : q <= 23'h250c22;
			12'd91   : q <= 23'h350c21;
			12'd92   : q <= 23'h21844e;
			12'd93   : q <= 23'h258042;
			12'd94   : q <= 23'h23b027;
			12'd95   : q <= 23'h298822;
			12'd96   : q <= 23'h241464;
			12'd97   : q <= 23'h354822;
			12'd98   : q <= 23'h34c822;
			12'd99   : q <= 23'h321d82;
			12'd100  : q <= 23'h31b842; 
			12'd101  : q <= 23'h353044; 
			12'd102  : q <= 23'h344822; 
			12'd103  : q <= 23'h358042; 
			12'd104  : q <= 23'h32b121; 
			12'd105  : q <= 23'h358042; 
			12'd106  : q <= 23'h3384c5; 
			12'd107  : q <= 23'h250042; 
			12'd108  : q <= 23'h31b421; 
			12'd109  : q <= 23'h343ca1; 
			12'd110  : q <= 23'h2290a6; 
			12'd111  : q <= 23'h34a924; 
			12'd112  : q <= 23'h2108c7; 
			12'd113  : q <= 23'h341c82; 
			12'd114  : q <= 23'h2398c2; 
			12'd115  : q <= 23'h222564; 
			12'd116  : q <= 23'h21b202; 
			12'd117  : q <= 23'h200601; 
			12'd118  : q <= 23'h349442; 
			12'd119  : q <= 23'h218865; 
			12'd120  : q <= 23'h352905; 
			12'd121  : q <= 23'h21b883; 
			12'd122  : q <= 23'h270c41; 
			12'd123  : q <= 23'h20b4e3; 
			12'd124  : q <= 23'h279043; 
			12'd125  : q <= 23'h2124e3; 
			12'd126  : q <= 23'h22a542; 
			12'd127  : q <= 23'h232484; 
			12'd128  : q <= 23'h270861; 
			12'd129  : q <= 23'h219042; 
			12'd130  : q <= 23'h25b844; 
			12'd131  : q <= 23'h3004a1; 
			12'd132  : q <= 23'h259524; 
			12'd133  : q <= 23'h232423; 
			12'd134  : q <= 23'h398821; 
			12'd135  : q <= 23'h349846; 
			12'd136  : q <= 23'h398821; 
			12'd137  : q <= 23'h31b841; 
			12'd138  : q <= 23'h261086; 
			12'd139  : q <= 23'h338843; 
			12'd140  : q <= 23'h231925; 
			12'd141  : q <= 23'h31104c; 
			12'd142  : q <= 23'h37b841; 
			12'd143  : q <= 23'h33bca1; 
			12'd144  : q <= 23'h37b861; 
			12'd145  : q <= 23'h333d01; 
			12'd146  : q <= 23'h37b861; 
			12'd147  : q <= 23'h313861; 
			12'd148  : q <= 23'h251cc6; 
			12'd149  : q <= 23'h251c26; 
			12'd150  : q <= 23'h2428a1; 
			12'd151  : q <= 23'h349824; 
			12'd152  : q <= 23'h24a844; 
			12'd153  : q <= 23'h341c26; 
			12'd154  : q <= 23'h360c23; 
			12'd155  : q <= 23'h339041; 
			12'd156  : q <= 23'h329d41; 
			12'd157  : q <= 23'h3398c3; 
			12'd158  : q <= 23'h349c61; 
			12'd159  : q <= 23'h213204; 
			12'd160  : q <= 23'h272443; 
			12'd161  : q <= 23'h30a8c5; 
			12'd162  : q <= 23'h350cc3; 
			12'd163  : q <= 23'h2334e7; 
			12'd164  : q <= 23'h36a462; 
			12'd165  : q <= 23'h3320a4; 
			12'd166  : q <= 23'h259c65; 
			12'd167  : q <= 23'h31a482; 
			12'd168  : q <= 23'h378c4a; 
			12'd169  : q <= 23'h229c85; 
			12'd170  : q <= 23'h2510c6; 
			12'd171  : q <= 23'h319049; 
			12'd172  : q <= 23'h258c25; 
			12'd173  : q <= 23'h240c25; 
			12'd174  : q <= 23'h353c41; 
			12'd175  : q <= 23'h243062; 
			12'd176  : q <= 23'h34bc41; 
			12'd177  : q <= 23'h223983; 
			12'd178  : q <= 23'h35b8a3; 
			12'd179  : q <= 23'h234061; 
			12'd180  : q <= 23'h360025; 
			12'd181  : q <= 23'h241467; 
			12'd182  : q <= 23'h368c23; 
			12'd183  : q <= 23'h218844; 
			12'd184  : q <= 23'h36b882; 
			12'd185  : q <= 23'h31b882; 
			12'd186  : q <= 23'h26b462; 
			12'd187  : q <= 23'h321481; 
			12'd188  : q <= 23'h23a564; 
			12'd189  : q <= 23'h342024; 
			12'd190  : q <= 23'h358441; 
			12'd191  : q <= 23'h329861; 
			12'd192  : q <= 23'h252543; 
			12'd193  : q <= 23'h349825; 
			12'd194  : q <= 23'h358421; 
			12'd195  : q <= 23'h220c81; 
			12'd196  : q <= 23'h361c81; 
			12'd197  : q <= 23'h338044; 
			12'd198  : q <= 23'h351c28; 
			12'd199  : q <= 23'h251c22; 
			12'd200  : q <= 23'h269ce2; 
			12'd201  : q <= 23'h301c62; 
			12'd202  : q <= 23'h26b462; 
			12'd203  : q <= 23'h223462; 
			12'd204  : q <= 23'h25a4c4; 
			12'd205  : q <= 23'h34b421; 
			12'd206  : q <= 23'h254442; 
			12'd207  : q <= 23'h349c41; 
			12'd208  : q <= 23'h278c63; 
			12'd209  : q <= 23'h301942; 
			12'd210  : q <= 23'h260c87; 
			12'd211  : q <= 23'h3224e5; 
			12'd212  : q <= 23'h278864; 
			12'd213  : q <= 23'h210864; 
			12'd214  : q <= 23'h3434c7; 
			12'd215  : q <= 23'h220c87; 
			12'd216  : q <= 23'h390c42; 
			12'd217  : q <= 23'h34b041; 
			12'd218  : q <= 23'h390c42; 
			12'd219  : q <= 23'h300c42; 
			12'd220  : q <= 23'h309e42; 
			12'd221  : q <= 23'h218867; 
			12'd222  : q <= 23'h23a8c7; 
			12'd223  : q <= 23'h21b1a5; 
			12'd224  : q <= 23'h25c041; 
			12'd225  : q <= 23'h212d02; 
			12'd226  : q <= 23'h281c62; 
			12'd227  : q <= 23'h333463; 
			12'd228  : q <= 23'h272423; 
			12'd229  : q <= 23'h23a841; 
			12'd230  : q <= 23'h3420a5; 
			12'd231  : q <= 23'h20a0a2; 
			12'd232  : q <= 23'h318e22; 
			12'd233  : q <= 23'h251c82; 
			12'd234  : q <= 23'h351c22; 
			12'd235  : q <= 23'h349c22; 
			12'd236  : q <= 23'h242881; 
			12'd237  : q <= 23'h342481; 
			12'd238  : q <= 23'h249464; 
			12'd239  : q <= 23'h343881; 
			12'd240  : q <= 23'h251cc3; 
			12'd241  : q <= 23'h343c81; 
			12'd242  : q <= 23'h34a061; 
			12'd243  : q <= 23'h341028; 
			12'd244  : q <= 23'h358026; 
			12'd245  : q <= 23'h240c48; 
			12'd246  : q <= 23'h270c6d; 
			12'd247  : q <= 23'h244063; 
			12'd248  : q <= 23'h270c6d; 
			12'd249  : q <= 23'h201ca2; 
			12'd250  : q <= 23'h270c6d; 
			12'd251  : q <= 23'h218c6d; 
			12'd252  : q <= 23'h248441; 
			12'd253  : q <= 23'h248021; 
			12'd254  : q <= 23'h264042; 
			12'd255  : q <= 23'h251823; 
			12'd256  : q <= 23'h341482; 
			12'd257  : q <= 23'h349c25; 
			12'd258  : q <= 23'h331902; 
			12'd259  : q <= 23'h24ac46; 
			12'd260  : q <= 23'h2228c4; 
			12'd261  : q <= 23'h260885; 
			12'd262  : q <= 23'h302641; 
			12'd263  : q <= 23'h244084; 
			12'd264  : q <= 23'h220885; 
			12'd265  : q <= 23'h26b462; 
			12'd266  : q <= 23'h33ac41; 
			12'd267  : q <= 23'h360c21; 
			12'd268  : q <= 23'h33b8a1; 
			12'd269  : q <= 23'h25b8e3; 
			12'd270  : q <= 23'h2138e3; 
			12'd271  : q <= 23'h364042; 
			12'd272  : q <= 23'h343c61; 
			12'd273  : q <= 23'h360025; 
			12'd274  : q <= 23'h240449; 
			12'd275  : q <= 23'h360c41; 
			12'd276  : q <= 23'h242862; 
			12'd277  : q <= 23'h243481; 
			12'd278  : q <= 23'h22cc81; 
			12'd279  : q <= 23'h310e42; 
			12'd280  : q <= 23'h338022; 
			12'd281  : q <= 23'h282061; 
			12'd282  : q <= 23'h233463; 
			12'd283  : q <= 23'h253542; 
			12'd284  : q <= 23'h349c45; 
			12'd285  : q <= 23'h258441; 
			12'd286  : q <= 23'h20a061; 
			12'd287  : q <= 23'h250941; 
			12'd288  : q <= 23'h33bca1; 
			12'd289  : q <= 23'h253463; 
			12'd290  : q <= 23'h34b441; 
			12'd291  : q <= 23'h383422; 
			12'd292  : q <= 23'h31b422; 
			12'd293  : q <= 23'h2590e6; 
			12'd294  : q <= 23'h329461; 
			12'd295  : q <= 23'h368c23; 
			12'd296  : q <= 23'h331d01; 
			12'd297  : q <= 23'h368c23; 
			12'd298  : q <= 23'h218445; 
			12'd299  : q <= 23'h229ca2; 
			12'd300  : q <= 23'h349c23; 
			12'd301  : q <= 23'h37b441; 
			12'd302  : q <= 23'h342024; 
			12'd303  : q <= 23'h26a826; 
			12'd304  : q <= 23'h2214c6; 
			12'd305  : q <= 23'h33bce1; 
			12'd306  : q <= 23'h31b441; 
			12'd307  : q <= 23'h2508e1; 
			12'd308  : q <= 23'h30842a; 
			12'd309  : q <= 23'h358045; 
			12'd310  : q <= 23'h241c62; 
			12'd311  : q <= 23'h2398c5; 
			12'd312  : q <= 23'h3384c3; 
			12'd313  : q <= 23'h381462; 
			12'd314  : q <= 23'h2318e3; 
			12'd315  : q <= 23'h341c82; 
			12'd316  : q <= 23'h202625; 
			12'd317  : q <= 23'h21b1e8; 
			12'd318  : q <= 23'h23c4c2; 
			12'd319  : q <= 23'h278849; 
			12'd320  : q <= 23'h211061; 
			12'd321  : q <= 23'h36a4e3; 
			12'd322  : q <= 23'h343081; 
			12'd323  : q <= 23'h250943; 
			12'd324  : q <= 23'h218865; 
			12'd325  : q <= 23'h26b062; 
			12'd326  : q <= 23'h223062; 
			12'd327  : q <= 23'h349443; 
			12'd328  : q <= 23'h23a8c4; 
			12'd329  : q <= 23'h203a83; 
			12'd330  : q <= 23'h223443; 
			12'd331  : q <= 23'h250086; 
			12'd332  : q <= 23'h2105e1; 
			12'd333  : q <= 23'h34b441; 
			12'd334  : q <= 23'h21b421; 
			12'd335  : q <= 23'h34b041; 
			12'd336  : q <= 23'h340c21; 
			12'd337  : q <= 23'h38a462; 
			12'd338  : q <= 23'h340822; 
			12'd339  : q <= 23'h3594a1; 
			12'd340  : q <= 23'h3214a1; 
			12'd341  : q <= 23'h299021; 
			12'd342  : q <= 23'h329881; 
			12'd343  : q <= 23'h38a462; 
			12'd344  : q <= 23'h302462; 
			12'd345  : q <= 23'h3714c3; 
			12'd346  : q <= 23'h3018a2; 
			12'd347  : q <= 23'h361442; 
			12'd348  : q <= 23'h331442; 
			12'd349  : q <= 23'h340c82; 
			12'd350  : q <= 23'h301062; 
			12'd351  : q <= 23'h331d01; 
			12'd352  : q <= 23'h3010a3; 
			12'd353  : q <= 23'h28004f; 
			12'd354  : q <= 23'h20ac61; 
			12'd355  : q <= 23'h272425; 
			12'd356  : q <= 23'h21044c; 
			12'd357  : q <= 23'h25ac42; 
			12'd358  : q <= 23'h23ac42; 
			12'd359  : q <= 23'h3420a5; 
			12'd360  : q <= 23'h21806a; 
			12'd361  : q <= 23'h361022; 
			12'd362  : q <= 23'h244064; 
			12'd363  : q <= 23'h343ca1; 
			12'd364  : q <= 23'h33bc81; 
			12'd365  : q <= 23'h361022; 
			12'd366  : q <= 23'h21bce2; 
			12'd367  : q <= 23'h250902; 
			12'd368  : q <= 23'h21a06c; 
			12'd369  : q <= 23'h229ca2; 
			12'd370  : q <= 23'h251c25; 
			12'd371  : q <= 23'h281c62; 
			12'd372  : q <= 23'h203901; 
			12'd373  : q <= 23'h281c62; 
			12'd374  : q <= 23'h209c62; 
			12'd375  : q <= 23'h263026; 
			12'd376  : q <= 23'h251426; 
			12'd377  : q <= 23'h373441; 
			12'd378  : q <= 23'h323441; 
			12'd379  : q <= 23'h343481; 
			12'd380  : q <= 23'h228822; 
			12'd381  : q <= 23'h329961; 
			12'd382  : q <= 23'h23b086; 
			12'd383  : q <= 23'h263485; 
			12'd384  : q <= 23'h23b026; 
			12'd385  : q <= 23'h220863; 
			12'd386  : q <= 23'h261465; 
			12'd387  : q <= 23'h229486; 
			12'd388  : q <= 23'h302682; 
			12'd389  : q <= 23'h220c41; 
			12'd390  : q <= 23'h344882; 
			12'd391  : q <= 23'h23b088; 
			12'd392  : q <= 23'h23a8e4; 
			12'd393  : q <= 23'h338c21; 
			12'd394  : q <= 23'h25c442; 
			12'd395  : q <= 23'h21a484; 
			12'd396  : q <= 23'h239cc6; 
			12'd397  : q <= 23'h331842; 
			12'd398  : q <= 23'h381882; 
			12'd399  : q <= 23'h2190a1; 
			12'd400  : q <= 23'h34b041; 
			12'd401  : q <= 23'h214481; 
			12'd402  : q <= 23'h253463; 
			12'd403  : q <= 23'h340024; 
			12'd404  : q <= 23'h344081; 
			12'd405  : q <= 23'h301882; 
			12'd406  : q <= 23'h349883; 
			12'd407  : q <= 23'h34984e; 
			12'd408  : q <= 23'h351c23; 
			12'd409  : q <= 23'h233842; 
			12'd410  : q <= 23'h3538e2; 
			12'd411  : q <= 23'h2085e1; 
			12'd412  : q <= 23'h270066; 
			12'd413  : q <= 23'h330c21; 
			12'd414  : q <= 23'h270066; 
			12'd415  : q <= 23'h202285; 
			12'd416  : q <= 23'h270066; 
			12'd417  : q <= 23'h218066; 
			12'd418  : q <= 23'h29c021; 
			12'd419  : q <= 23'h210848; 
			12'd420  : q <= 23'h258522; 
			12'd421  : q <= 23'h243421; 
			12'd422  : q <= 23'h2508a3; 
			12'd423  : q <= 23'h251c24; 
			12'd424  : q <= 23'h351c23; 
			12'd425  : q <= 23'h341488; 
			12'd426  : q <= 23'h37c081; 
			12'd427  : q <= 23'h34c821; 
			12'd428  : q <= 23'h34b881; 
			12'd429  : q <= 23'h33b881; 
			12'd430  : q <= 23'h29c021; 
			12'd431  : q <= 23'h204502; 
			12'd432  : q <= 23'h358c44; 
			12'd433  : q <= 23'h343c81; 
			12'd434  : q <= 23'h31c1c2; 
			12'd435  : q <= 23'h2318c3; 
			12'd436  : q <= 23'h22b943; 
			12'd437  : q <= 23'h322824; 
			12'd438  : q <= 23'h26a422; 
			12'd439  : q <= 23'h338c44; 
			12'd440  : q <= 23'h351c23; 
			12'd441  : q <= 23'h313441; 
			12'd442  : q <= 23'h34b064; 
			12'd443  : q <= 23'h21b843; 
			12'd444  : q <= 23'h284041; 
			12'd445  : q <= 23'h214041; 
			12'd446  : q <= 23'h343481; 
			12'd447  : q <= 23'h251d41; 
			12'd448  : q <= 23'h239883; 
			12'd449  : q <= 23'h249c82; 
			12'd450  : q <= 23'h351c25; 
			12'd451  : q <= 23'h349c25; 
			12'd452  : q <= 23'h360425; 
			12'd453  : q <= 23'h338826; 
			12'd454  : q <= 23'h273865; 
			12'd455  : q <= 23'h24a441; 
			12'd456  : q <= 23'h352021; 
			12'd457  : q <= 23'h231821; 
			12'd458  : q <= 23'h25ad22; 
			12'd459  : q <= 23'h231821; 
			12'd460  : q <= 23'h204281; 
			12'd461  : q <= 23'h323c41; 
			12'd462  : q <= 23'h343c81; 
			12'd463  : q <= 23'h342041; 
			12'd464  : q <= 23'h34ac41; 
			12'd465  : q <= 23'h229942; 
			12'd466  : q <= 23'h261c62; 
			12'd467  : q <= 23'h322462; 
			12'd468  : q <= 23'h26bc42; 
			12'd469  : q <= 23'h23a481; 
			12'd470  : q <= 23'h268443; 
			12'd471  : q <= 23'h22bc42; 
			12'd472  : q <= 23'h249447; 
			12'd473  : q <= 23'h249883; 
			12'd474  : q <= 23'h24a841; 
			12'd475  : q <= 23'h33c0a1; 
			12'd476  : q <= 23'h25a843; 
			12'd477  : q <= 23'h233905; 
			12'd478  : q <= 23'h252c62; 
			12'd479  : q <= 23'h23ac62; 
			12'd480  : q <= 23'h258c81; 
			12'd481  : q <= 23'h338c22; 
			12'd482  : q <= 23'h271465; 
			12'd483  : q <= 23'h23ac46; 
			12'd484  : q <= 23'h343081; 
			12'd485  : q <= 23'h228423; 
			12'd486  : q <= 23'h391442; 
			12'd487  : q <= 23'h301442; 
			12'd488  : q <= 23'h34b441; 
			12'd489  : q <= 23'h33b881; 
			12'd490  : q <= 23'h390842; 
			12'd491  : q <= 23'h300842; 
			12'd492  : q <= 23'h343cc1; 
			12'd493  : q <= 23'h241024; 
			12'd494  : q <= 23'h341c82; 
			12'd495  : q <= 23'h239022; 
			12'd496  : q <= 23'h2538e2; 
			12'd497  : q <= 23'h233c61; 
			12'd498  : q <= 23'h2740c1; 
			12'd499  : q <= 23'h214184; 
			12'd500  : q <= 23'h23a0e1; 
			12'd501  : q <= 23'h200e41; 
			12'd502  : q <= 23'h249825; 
			12'd503  : q <= 23'h341428; 
			12'd504  : q <= 23'h351824; 
			12'd505  : q <= 23'h223861; 
			12'd506  : q <= 23'h359043; 
			12'd507  : q <= 23'h339043; 
			12'd508  : q <= 23'h2730a1; 
			12'd509  : q <= 23'h318849; 
			12'd510  : q <= 23'h27186d; 
			12'd511  : q <= 23'h2198e4; 
			12'd512  : q <= 23'h28004b; 
			12'd513  : q <= 23'h2190c6; 
			12'd514  : q <= 23'h3594a1; 
			12'd515  : q <= 23'h223081; 
			12'd516  : q <= 23'h251c22; 
			12'd517  : q <= 23'h249c22; 
			12'd518  : q <= 23'h354422; 
			12'd519  : q <= 23'h329c61; 
			12'd520  : q <= 23'h358023; 
			12'd521  : q <= 23'h229861; 
			12'd522  : q <= 23'h364481; 
			12'd523  : q <= 23'h21b461; 
			12'd524  : q <= 23'h24b461; 
			12'd525  : q <= 23'h20ad02; 
			12'd526  : q <= 23'h361461; 
			12'd527  : q <= 23'h3214a1; 
			12'd528  : q <= 23'h364481; 
			12'd529  : q <= 23'h329461; 
			12'd530  : q <= 23'h248441; 
			12'd531  : q <= 23'h242881; 
			12'd532  : q <= 23'h342481; 
			12'd533  : q <= 23'h313443; 
			12'd534  : q <= 23'h283c61; 
			12'd535  : q <= 23'h33c8c2; 
			12'd536  : q <= 23'h283c61; 
			12'd537  : q <= 23'h20bc61; 
			12'd538  : q <= 23'h33bcc1; 
			12'd539  : q <= 23'h32bd01; 
			12'd540  : q <= 23'h25184e; 
			12'd541  : q <= 23'h24184e; 
			12'd542  : q <= 23'h369841; 
			12'd543  : q <= 23'h34c041; 
			12'd544  : q <= 23'h34b461; 
			12'd545  : q <= 23'h340023; 
			12'd546  : q <= 23'h222609; 
			12'd547  : q <= 23'h20a207; 
			12'd548  : q <= 23'h3424a4; 
			12'd549  : q <= 23'h3334e1; 
			12'd550  : q <= 23'h374041; 
			12'd551  : q <= 23'h210d07; 
			12'd552  : q <= 23'h290849; 
			12'd553  : q <= 23'h324041; 
			12'd554  : q <= 23'h290849; 
			12'd555  : q <= 23'h308901; 
			12'd556  : q <= 23'h343081; 
			12'd557  : q <= 23'h32b8a3; 
			12'd558  : q <= 23'h28004b; 
			12'd559  : q <= 23'h348041; 
			12'd560  : q <= 23'h388c27; 
			12'd561  : q <= 23'h310c27; 
			12'd562  : q <= 23'h33b0c4; 
			12'd563  : q <= 23'h21004b; 
			12'd564  : q <= 23'h270074; 
			12'd565  : q <= 23'h201021; 
			12'd566  : q <= 23'h2514a4; 
			12'd567  : q <= 23'h221cc2; 
			12'd568  : q <= 23'h228464; 
			12'd569  : q <= 23'h261c62; 
			12'd570  : q <= 23'h22a443; 
			12'd571  : q <= 23'h264062; 
			12'd572  : q <= 23'h24a846; 
			12'd573  : q <= 23'h348452; 
			12'd574  : q <= 23'h343082; 
			12'd575  : q <= 23'h2424c1; 
			12'd576  : q <= 23'h348026; 
			12'd577  : q <= 23'h25cc61; 
			12'd578  : q <= 23'h208e22; 
			12'd579  : q <= 23'h25a04c; 
			12'd580  : q <= 23'h343c81; 
			12'd581  : q <= 23'h260c31; 
			12'd582  : q <= 23'h331c41; 
			12'd583  : q <= 23'h391041; 
			12'd584  : q <= 23'h241862; 
			12'd585  : q <= 23'h222985; 
			12'd586  : q <= 23'h23c842; 
			12'd587  : q <= 23'h389062; 
			12'd588  : q <= 23'h349c46; 
			12'd589  : q <= 23'h389062; 
			12'd590  : q <= 23'h348024; 
			12'd591  : q <= 23'h34bc41; 
			12'd592  : q <= 23'h3034c1; 
			12'd593  : q <= 23'h343c81; 
			12'd594  : q <= 23'h31b441; 
			12'd595  : q <= 23'h349887; 
			12'd596  : q <= 23'h301062; 
			12'd597  : q <= 23'h371c21; 
			12'd598  : q <= 23'h31802e; 
			12'd599  : q <= 23'h3640a2; 
			12'd600  : q <= 23'h3240a2; 
			12'd601  : q <= 23'h262821; 
			12'd602  : q <= 23'h33002e; 
			12'd603  : q <= 23'h354041; 
			12'd604  : q <= 23'h300c41; 
			12'd605  : q <= 23'h22b983; 
			12'd606  : q <= 23'h333863; 
			12'd607  : q <= 23'h262821; 
			12'd608  : q <= 23'h329c21; 
			12'd609  : q <= 23'h3229a1; 
			12'd610  : q <= 23'h331ca6; 
			12'd611  : q <= 23'h341486; 
			12'd612  : q <= 23'h342c81; 
			12'd613  : q <= 23'h37bc21; 
			12'd614  : q <= 23'h30b0a1; 
			12'd615  : q <= 23'h239ce6; 
			12'd616  : q <= 23'h200465; 
			12'd617  : q <= 23'h380881; 
			12'd618  : q <= 23'h329841; 
			12'd619  : q <= 23'h368825; 
			12'd620  : q <= 23'h301482; 
			12'd621  : q <= 23'h243481; 
			12'd622  : q <= 23'h34c821; 
			12'd623  : q <= 23'h262821; 
			12'd624  : q <= 23'h23a821; 
			12'd625  : q <= 23'h25b482; 
			12'd626  : q <= 23'h34b028; 
			12'd627  : q <= 23'h3684c1; 
			12'd628  : q <= 23'h34a024; 
			12'd629  : q <= 23'h251ca5; 
			12'd630  : q <= 23'h21c881; 
			12'd631  : q <= 23'h360848; 
			12'd632  : q <= 23'h330848; 
			12'd633  : q <= 23'h360027; 
			12'd634  : q <= 23'h242c21; 
			12'd635  : q <= 23'h37bc21; 
			12'd636  : q <= 23'h23bc21; 
			12'd637  : q <= 23'h37bc21; 
			12'd638  : q <= 23'h338027; 
			12'd639  : q <= 23'h290427; 
			12'd640  : q <= 23'h21290a; 
			12'd641  : q <= 23'h3189e2; 
			12'd642  : q <= 23'h221181; 
			12'd643  : q <= 23'h280045; 
			12'd644  : q <= 23'h340024; 
			12'd645  : q <= 23'h280045; 
			12'd646  : q <= 23'h319c4d; 
			12'd647  : q <= 23'h280045; 
			12'd648  : q <= 23'h210045; 
			12'd649  : q <= 23'h373862; 
			12'd650  : q <= 23'h31b862; 
			12'd651  : q <= 23'h380881; 
			12'd652  : q <= 23'h241c25; 
			12'd653  : q <= 23'h25b482; 
			12'd654  : q <= 23'h300881; 
			12'd655  : q <= 23'h369421; 
			12'd656  : q <= 23'h343c25; 
			12'd657  : q <= 23'h351c25; 
			12'd658  : q <= 23'h349c25; 
			12'd659  : q <= 23'h25184e; 
			12'd660  : q <= 23'h301ca2; 
			12'd661  : q <= 23'h249464; 
			12'd662  : q <= 23'h3300ca; 
			12'd663  : q <= 23'h25184e; 
			12'd664  : q <= 23'h24184e; 
			12'd665  : q <= 23'h369421; 
			12'd666  : q <= 23'h230423; 
			12'd667  : q <= 23'h298429; 
			12'd668  : q <= 23'h310881; 
			12'd669  : q <= 23'h298429; 
			12'd670  : q <= 23'h20b843; 
			12'd671  : q <= 23'h3534e2; 
			12'd672  : q <= 23'h202865; 
			12'd673  : q <= 23'h360024; 
			12'd674  : q <= 23'h22b4a3; 
			12'd675  : q <= 23'h272824; 
			12'd676  : q <= 23'h209d23; 
			12'd677  : q <= 23'h249c22; 
			12'd678  : q <= 23'h23a445; 
			12'd679  : q <= 23'h349843; 
			12'd680  : q <= 23'h3380c4; 
			12'd681  : q <= 23'h23c442; 
			12'd682  : q <= 23'h308e63; 
			12'd683  : q <= 23'h31a462; 
			12'd684  : q <= 23'h279c42; 
			12'd685  : q <= 23'h219c42; 
			12'd686  : q <= 23'h24a944; 
			12'd687  : q <= 23'h21b9c6; 
			12'd688  : q <= 23'h2594a6; 
			12'd689  : q <= 23'h34b041; 
			12'd690  : q <= 23'h249465; 
			12'd691  : q <= 23'h249842; 
			12'd692  : q <= 23'h249465; 
			12'd693  : q <= 23'h241465; 
			12'd694  : q <= 23'h368841; 
			12'd695  : q <= 23'h328841; 
			12'd696  : q <= 23'h369841; 
			12'd697  : q <= 23'h203022; 
			12'd698  : q <= 23'h369841; 
			12'd699  : q <= 23'h34c822; 
			12'd700  : q <= 23'h234121; 
			12'd701  : q <= 23'h343c81; 
			12'd702  : q <= 23'h291842; 
			12'd703  : q <= 23'h329841; 
			12'd704  : q <= 23'h27c461; 
			12'd705  : q <= 23'h300c63; 
			12'd706  : q <= 23'h34a061; 
			12'd707  : q <= 23'h342061; 
			12'd708  : q <= 23'h249426; 
			12'd709  : q <= 23'h349824; 
			12'd710  : q <= 23'h259886; 
			12'd711  : q <= 23'h229886; 
			12'd712  : q <= 23'h361461; 
			12'd713  : q <= 23'h214461; 
			12'd714  : q <= 23'h361461; 
			12'd715  : q <= 23'h3138c2; 
			12'd716  : q <= 23'h33b8c1; 
			12'd717  : q <= 23'h333cc1; 
			12'd718  : q <= 23'h3740a1; 
			12'd719  : q <= 23'h329461; 
			12'd720  : q <= 23'h3740a1; 
			12'd721  : q <= 23'h338c42; 
			12'd722  : q <= 23'h344081; 
			12'd723  : q <= 23'h30c0a1; 
			12'd724  : q <= 23'h253443; 
			12'd725  : q <= 23'h342023; 
			12'd726  : q <= 23'h2608a2; 
			12'd727  : q <= 23'h200941; 
			12'd728  : q <= 23'h3380c4; 
			12'd729  : q <= 23'h330c41; 
			12'd730  : q <= 23'h224da1; 
			12'd731  : q <= 23'h313062; 
			12'd732  : q <= 23'h28b064; 
			12'd733  : q <= 23'h2234a3; 
			12'd734  : q <= 23'h273421; 
			12'd735  : q <= 23'h343881; 
			12'd736  : q <= 23'h273441; 
			12'd737  : q <= 23'h223441; 
			12'd738  : q <= 23'h243521; 
			12'd739  : q <= 23'h34bc41; 
			12'd740  : q <= 23'h25b463; 
			12'd741  : q <= 23'h22b126; 
			12'd742  : q <= 23'h25b463; 
			12'd743  : q <= 23'h233463; 
			12'd744  : q <= 23'h329561; 
			12'd745  : q <= 23'h2398a5; 
			12'd746  : q <= 23'h212641; 
			12'd747  : q <= 23'h33c8a1; 
			12'd748  : q <= 23'h34a481; 
			12'd749  : q <= 23'h203863; 
			12'd750  : q <= 23'h34a481; 
			12'd751  : q <= 23'h33a481; 
			12'd752  : q <= 23'h272867; 
			12'd753  : q <= 23'h208601; 
			12'd754  : q <= 23'h353143; 
			12'd755  : q <= 23'h2284a2; 
			12'd756  : q <= 23'h389041; 
			12'd757  : q <= 23'h309041; 
			12'd758  : q <= 23'h351c26; 
			12'd759  : q <= 23'h241443; 
			12'd760  : q <= 23'h349446; 
			12'd761  : q <= 23'h2190c6; 
			12'd762  : q <= 23'h35884f; 
			12'd763  : q <= 23'h320851; 
			12'd764  : q <= 23'h272867; 
			12'd765  : q <= 23'h21a867; 
			12'd766  : q <= 23'h35884f; 
			12'd767  : q <= 23'h33884f; 
			12'd768  : q <= 23'h38ac62; 
			12'd769  : q <= 23'h341c46; 
			12'd770  : q <= 23'h252923; 
			12'd771  : q <= 23'h303143; 
			12'd772  : q <= 23'h344081; 
			12'd773  : q <= 23'h22b862; 
			12'd774  : q <= 23'h21a606; 
			12'd775  : q <= 23'h2084c6; 
			12'd776  : q <= 23'h259022; 
			12'd777  : q <= 23'h2024a1; 
			12'd778  : q <= 23'h34b061; 
			12'd779  : q <= 23'h21b521; 
			12'd780  : q <= 23'h24a841; 
			12'd781  : q <= 23'h3199a2; 
			12'd782  : q <= 23'h261c62; 
			12'd783  : q <= 23'h220068; 
			12'd784  : q <= 23'h24ac46; 
			12'd785  : q <= 23'h222465; 
			12'd786  : q <= 23'h334901; 
			12'd787  : q <= 23'h301d42; 
			12'd788  : q <= 23'h268c61; 
			12'd789  : q <= 23'h249445; 
			12'd790  : q <= 23'h364062; 
			12'd791  : q <= 23'h20b101; 
			12'd792  : q <= 23'h33b8c1; 
			12'd793  : q <= 23'h301c62; 
			12'd794  : q <= 23'h268c61; 
			12'd795  : q <= 23'h223843; 
			12'd796  : q <= 23'h268c61; 
			12'd797  : q <= 23'h341884; 
			12'd798  : q <= 23'h288064; 
			12'd799  : q <= 23'h344422; 
			12'd800  : q <= 23'h243481; 
			12'd801  : q <= 23'h230086; 
			12'd802  : q <= 23'h278025; 
			12'd803  : q <= 23'h228c83; 
			12'd804  : q <= 23'h288065; 
			12'd805  : q <= 23'h24bc21; 
			12'd806  : q <= 23'h37ac81; 
			12'd807  : q <= 23'h343c41; 
			12'd808  : q <= 23'h2534e2; 
			12'd809  : q <= 23'h30ac81; 
			12'd810  : q <= 23'h35ac41; 
			12'd811  : q <= 23'h33ac41; 
			12'd812  : q <= 23'h31aa05; 
			12'd813  : q <= 23'h243042; 
			12'd814  : q <= 23'h2510c5; 
			12'd815  : q <= 23'h349824; 
			12'd816  : q <= 23'h253044; 
			12'd817  : q <= 23'h343c81; 
			12'd818  : q <= 23'h368822; 
			12'd819  : q <= 23'h244061; 
			12'd820  : q <= 23'h34806e; 
			12'd821  : q <= 23'h251823; 
			12'd822  : q <= 23'h352441; 
			12'd823  : q <= 23'h302c82; 
			12'd824  : q <= 23'h230501; 
			12'd825  : q <= 23'h333ce1; 
			12'd826  : q <= 23'h343503; 
			12'd827  : q <= 23'h330822; 
			12'd828  : q <= 23'h288464; 
			12'd829  : q <= 23'h200464; 
			12'd830  : q <= 23'h250923; 
			12'd831  : q <= 23'h250c21; 
			12'd832  : q <= 23'h278843; 
			12'd833  : q <= 23'h329461; 
			12'd834  : q <= 23'h369821; 
			12'd835  : q <= 23'h3144a1; 
			12'd836  : q <= 23'h278843; 
			12'd837  : q <= 23'h218843; 
			12'd838  : q <= 23'h269821; 
			12'd839  : q <= 23'h229841; 
			12'd840  : q <= 23'h26a422; 
			12'd841  : q <= 23'h232422; 
			12'd842  : q <= 23'h26c861; 
			12'd843  : q <= 23'h234042; 
			12'd844  : q <= 23'h34c441; 
			12'd845  : q <= 23'h303d22; 
			12'd846  : q <= 23'h24c443; 
			12'd847  : q <= 23'h34c041; 
			12'd848  : q <= 23'h30b242; 
			12'd849  : q <= 23'h243081; 
			12'd850  : q <= 23'h23a8c1; 
			12'd851  : q <= 23'h342441; 
			12'd852  : q <= 23'h391424; 
			12'd853  : q <= 23'h33ccc1; 
			12'd854  : q <= 23'h350022; 
			12'd855  : q <= 23'h30a822; 
			12'd856  : q <= 23'h264483; 
			12'd857  : q <= 23'h309424; 
			12'd858  : q <= 23'h34a041; 
			12'd859  : q <= 23'h23ac21; 
			12'd860  : q <= 23'h258c25; 
			12'd861  : q <= 23'h240c25; 
			12'd862  : q <= 23'h37b841; 
			12'd863  : q <= 23'h329c41; 
			12'd864  : q <= 23'h34cca1; 
			12'd865  : q <= 23'h334ca1; 
			12'd866  : q <= 23'h37b841; 
			12'd867  : q <= 23'h23804f; 
			12'd868  : q <= 23'h249825; 
			12'd869  : q <= 23'h251427; 
			12'd870  : q <= 23'h383061; 
			12'd871  : q <= 23'h30b061; 
			12'd872  : q <= 23'h331d01; 
			12'd873  : q <= 23'h2040c1; 
			12'd874  : q <= 23'h3380c6; 
			12'd875  : q <= 23'h338024; 
			12'd876  : q <= 23'h282845; 
			12'd877  : q <= 23'h320822; 
			12'd878  : q <= 23'h258c41; 
			12'd879  : q <= 23'h212845; 
			12'd880  : q <= 23'h253543; 
			12'd881  : q <= 23'h20942f; 
			12'd882  : q <= 23'h251d22; 
			12'd883  : q <= 23'h208031; 
			12'd884  : q <= 23'h251903; 
			12'd885  : q <= 23'h343c21; 
			12'd886  : q <= 23'h244081; 
			12'd887  : q <= 23'h228881; 
			12'd888  : q <= 23'h233903; 
			12'd889  : q <= 23'h24b841; 
			12'd890  : q <= 23'h391842; 
			12'd891  : q <= 23'h24b441; 
			12'd892  : q <= 23'h391842; 
			12'd893  : q <= 23'h34b821; 
			12'd894  : q <= 23'h391842; 
			12'd895  : q <= 23'h301842; 
			12'd896  : q <= 23'h34b461; 
			12'd897  : q <= 23'h31b841; 
			12'd898  : q <= 23'h36b881; 
			12'd899  : q <= 23'h329461; 
			12'd900  : q <= 23'h329142; 
			12'd901  : q <= 23'h31b881; 
			12'd902  : q <= 23'h341ca5; 
			12'd903  : q <= 23'h339c82; 
			12'd904  : q <= 23'h358c29; 
			12'd905  : q <= 23'h251846; 
			12'd906  : q <= 23'h34a081; 
			12'd907  : q <= 23'h212449; 
			12'd908  : q <= 23'h353425; 
			12'd909  : q <= 23'h349c43; 
			12'd910  : q <= 23'h351c25; 
			12'd911  : q <= 23'h249c82; 
			12'd912  : q <= 23'h34a482; 
			12'd913  : q <= 23'h2518a3; 
			12'd914  : q <= 23'h35b021; 
			12'd915  : q <= 23'h301965; 
			12'd916  : q <= 23'h3380c6; 
			12'd917  : q <= 23'h349c41; 
			12'd918  : q <= 23'h22c062; 
			12'd919  : q <= 23'h232524; 
			12'd920  : q <= 23'h22b443; 
			12'd921  : q <= 23'h259885; 
			12'd922  : q <= 23'h229885; 
			12'd923  : q <= 23'h249841; 
			12'd924  : q <= 23'h22b501; 
			12'd925  : q <= 23'h250d01; 
			12'd926  : q <= 23'h220025; 
			12'd927  : q <= 23'h24ac41; 
			12'd928  : q <= 23'h3125e1; 
			12'd929  : q <= 23'h343881; 
			12'd930  : q <= 23'h340822; 
			12'd931  : q <= 23'h33b8c1; 
			12'd932  : q <= 23'h24a841; 
			12'd933  : q <= 23'h389062; 
			12'd934  : q <= 23'h311424; 
			12'd935  : q <= 23'h372882; 
			12'd936  : q <= 23'h311028; 
			12'd937  : q <= 23'h244083; 
			12'd938  : q <= 23'h21bc41; 
			12'd939  : q <= 23'h372882; 
			12'd940  : q <= 23'h312882; 
			12'd941  : q <= 23'h254423; 
			12'd942  : q <= 23'h341426; 
			12'd943  : q <= 23'h260823; 
			12'd944  : q <= 23'h341845; 
			12'd945  : q <= 23'h388c62; 
			12'd946  : q <= 23'h349c25; 
			12'd947  : q <= 23'h354822; 
			12'd948  : q <= 23'h34c822; 
			12'd949  : q <= 23'h2610a1; 
			12'd950  : q <= 23'h239ca6; 
			12'd951  : q <= 23'h3380c4; 
			12'd952  : q <= 23'h220c41; 
			12'd953  : q <= 23'h26b841; 
			12'd954  : q <= 23'h301062; 
			12'd955  : q <= 23'h34a041; 
			12'd956  : q <= 23'h329821; 
			12'd957  : q <= 23'h252861; 
			12'd958  : q <= 23'h23a861; 
			12'd959  : q <= 23'h34c861; 
			12'd960  : q <= 23'h323c21; 
			12'd961  : q <= 23'h361861; 
			12'd962  : q <= 23'h321981; 
			12'd963  : q <= 23'h34a441; 
			12'd964  : q <= 23'h32a423; 
			12'd965  : q <= 23'h348071; 
			12'd966  : q <= 23'h34b421; 
			12'd967  : q <= 23'h34a845; 
			12'd968  : q <= 23'h343c41; 
			12'd969  : q <= 23'h353c21; 
			12'd970  : q <= 23'h348445; 
			12'd971  : q <= 23'h200142; 
			12'd972  : q <= 23'h3138a1; 
			12'd973  : q <= 23'h34b041; 
			12'd974  : q <= 23'h312925; 
			12'd975  : q <= 23'h2580c5; 
			12'd976  : q <= 23'h230423; 
			12'd977  : q <= 23'h361c41; 
			12'd978  : q <= 23'h218425; 
			12'd979  : q <= 23'h269c21; 
			12'd980  : q <= 23'h323c82; 
			12'd981  : q <= 23'h269c21; 
			12'd982  : q <= 23'h231c21; 
			12'd983  : q <= 23'h25b122; 
			12'd984  : q <= 23'h229c21; 
			12'd985  : q <= 23'h281081; 
			12'd986  : q <= 23'h200829; 
			12'd987  : q <= 23'h250922; 
			12'd988  : q <= 23'h34bc21; 
			12'd989  : q <= 23'h25b122; 
			12'd990  : q <= 23'h203122; 
			12'd991  : q <= 23'h3594a1; 
			12'd992  : q <= 23'h3314e1; 
			12'd993  : q <= 23'h36c861; 
			12'd994  : q <= 23'h348424; 
			12'd995  : q <= 23'h259024; 
			12'd996  : q <= 23'h31c463; 
			12'd997  : q <= 23'h260024; 
			12'd998  : q <= 23'h202066; 
			12'd999  : q <= 23'h253486; 
			12'd1000 : q <= 23'h22a907; 
			12'd1001 : q <= 23'h272861; 
			12'd1002 : q <= 23'h201942; 
			12'd1003 : q <= 23'h2510a4; 
			12'd1004 : q <= 23'h240444; 
			12'd1005 : q <= 23'h35ac41; 
			12'd1006 : q <= 23'h34a424; 
			12'd1007 : q <= 23'h391842; 
			12'd1008 : q <= 23'h34a024; 
			12'd1009 : q <= 23'h3389a1; 
			12'd1010 : q <= 23'h34b441; 
			12'd1011 : q <= 23'h363462; 
			12'd1012 : q <= 23'h33ac41; 
			12'd1013 : q <= 23'h251125; 
			12'd1014 : q <= 23'h342483; 
			12'd1015 : q <= 23'h341c81; 
			12'd1016 : q <= 23'h349c23; 
			12'd1017 : q <= 23'h374081; 
			12'd1018 : q <= 23'h33282a; 
			12'd1019 : q <= 23'h344081; 
			12'd1020 : q <= 23'h302822; 
			12'd1021 : q <= 23'h354021; 
			12'd1022 : q <= 23'h314081; 
			12'd1023 : q <= 23'h298c24; 
			12'd1024 : q <= 23'h200c24; 
			12'd1025 : q <= 23'h251ce5; 
			12'd1026 : q <= 23'h302261; 
			12'd1027 : q <= 23'h361c61; 
			12'd1028 : q <= 23'h301c21; 
			12'd1029 : q <= 23'h361c61; 
			12'd1030 : q <= 23'h329c61; 
			12'd1031 : q <= 23'h240c81; 
			12'd1032 : q <= 23'h240c4c; 
			12'd1033 : q <= 23'h369c41; 
			12'd1034 : q <= 23'h203282; 
			12'd1035 : q <= 23'h211e27; 
			12'd1036 : q <= 23'h200065; 
			12'd1037 : q <= 23'h271864; 
			12'd1038 : q <= 23'h219864; 
			12'd1039 : q <= 23'h268ce1; 
			12'd1040 : q <= 23'h200ce1; 
			12'd1041 : q <= 23'h26ace1; 
			12'd1042 : q <= 23'h241421; 
			12'd1043 : q <= 23'h26a423; 
			12'd1044 : q <= 23'h31042c; 
			12'd1045 : q <= 23'h389421; 
			12'd1046 : q <= 23'h311421; 
			12'd1047 : q <= 23'h371821; 
			12'd1048 : q <= 23'h33c441; 
			12'd1049 : q <= 23'h253443; 
			12'd1050 : q <= 23'h329821; 
			12'd1051 : q <= 23'h280054; 
			12'd1052 : q <= 23'h228423; 
			12'd1053 : q <= 23'h229942; 
			12'd1054 : q <= 23'h27884c; 
			12'd1055 : q <= 23'h23b086; 
			12'd1056 : q <= 23'h272424; 
			12'd1057 : q <= 23'h2090e5; 
			12'd1058 : q <= 23'h271867; 
			12'd1059 : q <= 23'h219867; 
			12'd1060 : q <= 23'h34a4a2; 
			12'd1061 : q <= 23'h33bcc1; 
			12'd1062 : q <= 23'h268ce2; 
			12'd1063 : q <= 23'h3324a2; 
			12'd1064 : q <= 23'h333903; 
			12'd1065 : q <= 23'h341028; 
			12'd1066 : q <= 23'h272443; 
			12'd1067 : q <= 23'h229c62; 
			12'd1068 : q <= 23'h3384d3; 
			12'd1069 : q <= 23'h220865; 
			12'd1070 : q <= 23'h2648c1; 
			12'd1071 : q <= 23'h2148c1; 
			12'd1072 : q <= 23'h389462; 
			12'd1073 : q <= 23'h344861; 
			12'd1074 : q <= 23'h254043; 
			12'd1075 : q <= 23'h33b8c1; 
			12'd1076 : q <= 23'h389462; 
			12'd1077 : q <= 23'h343841; 
			12'd1078 : q <= 23'h358c42; 
			12'd1079 : q <= 23'h301462; 
			12'd1080 : q <= 23'h341c82; 
			12'd1081 : q <= 23'h229861; 
			12'd1082 : q <= 23'h358424; 
			12'd1083 : q <= 23'h3094a3; 
			12'd1084 : q <= 23'h369c41; 
			12'd1085 : q <= 23'h2398e3; 
			12'd1086 : q <= 23'h213e44; 
			12'd1087 : q <= 23'h329c41; 
			12'd1088 : q <= 23'h261841; 
			12'd1089 : q <= 23'h231841; 
			12'd1090 : q <= 23'h358424; 
			12'd1091 : q <= 23'h240427; 
			12'd1092 : q <= 23'h2225e7; 
			12'd1093 : q <= 23'h349c22; 
			12'd1094 : q <= 23'h258d22; 
			12'd1095 : q <= 23'h251c22; 
			12'd1096 : q <= 23'h26a423; 
			12'd1097 : q <= 23'h338842; 
			12'd1098 : q <= 23'h249427; 
			12'd1099 : q <= 23'h232423; 
			12'd1100 : q <= 23'h2325c9; 
			12'd1101 : q <= 23'h3144c1; 
			12'd1102 : q <= 23'h351c26; 
			12'd1103 : q <= 23'h33a481; 
			12'd1104 : q <= 23'h33b4c1; 
			12'd1105 : q <= 23'h34b441; 
			12'd1106 : q <= 23'h34b042; 
			12'd1107 : q <= 23'h22b883; 
			12'd1108 : q <= 23'h25b4e1; 
			12'd1109 : q <= 23'h232883; 
			12'd1110 : q <= 23'h25b062; 
			12'd1111 : q <= 23'h34c441; 
			12'd1112 : q <= 23'h369823; 
			12'd1113 : q <= 23'h30bdc2; 
			12'd1114 : q <= 23'h26a423; 
			12'd1115 : q <= 23'h309028; 
			12'd1116 : q <= 23'h290032; 
			12'd1117 : q <= 23'h2110c1; 
			12'd1118 : q <= 23'h348902; 
			12'd1119 : q <= 23'h232423; 
			12'd1120 : q <= 23'h3724c1; 
			12'd1121 : q <= 23'h208032; 
			12'd1122 : q <= 23'h254921; 
			12'd1123 : q <= 23'h21c041; 
			12'd1124 : q <= 23'h343ca1; 
			12'd1125 : q <= 23'h343c41; 
			12'd1126 : q <= 23'h368c23; 
			12'd1127 : q <= 23'h349442; 
			12'd1128 : q <= 23'h2798a1; 
			12'd1129 : q <= 23'h2018a1; 
			12'd1130 : q <= 23'h28c423; 
			12'd1131 : q <= 23'h32a463; 
			12'd1132 : q <= 23'h368c23; 
			12'd1133 : q <= 23'h210052; 
			12'd1134 : q <= 23'h389c21; 
			12'd1135 : q <= 23'h214423; 
			12'd1136 : q <= 23'h29a421; 
			12'd1137 : q <= 23'h330c23; 
			12'd1138 : q <= 23'h34c441; 
			12'd1139 : q <= 23'h311c21; 
			12'd1140 : q <= 23'h281081; 
			12'd1141 : q <= 23'h201081; 
			12'd1142 : q <= 23'h214a42; 
			12'd1143 : q <= 23'h23c442; 
			12'd1144 : q <= 23'h3205c1; 
			12'd1145 : q <= 23'h210054; 
			12'd1146 : q <= 23'h271044; 
			12'd1147 : q <= 23'h231c21; 
			12'd1148 : q <= 23'h351c41; 
			12'd1149 : q <= 23'h242061; 
			12'd1150 : q <= 23'h2420c6; 
			12'd1151 : q <= 23'h321164; 
			12'd1152 : q <= 23'h38244b; 
			12'd1153 : q <= 23'h303c81; 
			12'd1154 : q <= 23'h34ac41; 
			12'd1155 : q <= 23'h22b061; 
			12'd1156 : q <= 23'h353c23; 
			12'd1157 : q <= 23'h34a024; 
			12'd1158 : q <= 23'h353c23; 
			12'd1159 : q <= 23'h341c22; 
			12'd1160 : q <= 23'h252902; 
			12'd1161 : q <= 23'h220c51; 
			12'd1162 : q <= 23'h27b427; 
			12'd1163 : q <= 23'h228861; 
			12'd1164 : q <= 23'h348884; 
			12'd1165 : q <= 23'h230086; 
			12'd1166 : q <= 23'h271c21; 
			12'd1167 : q <= 23'h303a82; 
			12'd1168 : q <= 23'h271c23; 
			12'd1169 : q <= 23'h31a06c; 
			12'd1170 : q <= 23'h218102; 
			12'd1171 : q <= 23'h334061; 
			12'd1172 : q <= 23'h3440c1; 
			12'd1173 : q <= 23'h303022; 
			12'd1174 : q <= 23'h352881; 
			12'd1175 : q <= 23'h34c041; 
			12'd1176 : q <= 23'h229ca1; 
			12'd1177 : q <= 23'h2500d3; 
			12'd1178 : q <= 23'h251943; 
			12'd1179 : q <= 23'h219821; 
			12'd1180 : q <= 23'h281821; 
			12'd1181 : q <= 23'h219821; 
			12'd1182 : q <= 23'h272826; 
			12'd1183 : q <= 23'h211505; 
			12'd1184 : q <= 23'h354422; 
			12'd1185 : q <= 23'h209441; 
			12'd1186 : q <= 23'h3500a5; 
			12'd1187 : q <= 23'h3280a5; 
			12'd1188 : q <= 23'h258831; 
			12'd1189 : q <= 23'h240831; 
			12'd1190 : q <= 23'h27ac29; 
			12'd1191 : q <= 23'h222c29; 
			12'd1192 : q <= 23'h22c0e4; 
			12'd1193 : q <= 23'h3390c1; 
			12'd1194 : q <= 23'h281c62; 
			12'd1195 : q <= 23'h34b044; 
			12'd1196 : q <= 23'h360cc2; 
			12'd1197 : q <= 23'h228863; 
			12'd1198 : q <= 23'h264062; 
			12'd1199 : q <= 23'h3388c3; 
			12'd1200 : q <= 23'h23a525; 
			12'd1201 : q <= 23'h23a444; 
			12'd1202 : q <= 23'h25b463; 
			12'd1203 : q <= 23'h33b0a1; 
			12'd1204 : q <= 23'h252c63; 
			12'd1205 : q <= 23'h300d43; 
			12'd1206 : q <= 23'h36c022; 
			12'd1207 : q <= 23'h301062; 
			12'd1208 : q <= 23'h343c81; 
			12'd1209 : q <= 23'h334022; 
			12'd1210 : q <= 23'h34c041; 
			12'd1211 : q <= 23'h339023; 
			12'd1212 : q <= 23'h348561; 
			12'd1213 : q <= 23'h301e81; 
			12'd1214 : q <= 23'h250821; 
			12'd1215 : q <= 23'h251826; 
			12'd1216 : q <= 23'h34a081; 
			12'd1217 : q <= 23'h33a081; 
			12'd1218 : q <= 23'h351c25; 
			12'd1219 : q <= 23'h232462; 
			12'd1220 : q <= 23'h362861; 
			12'd1221 : q <= 23'h348041; 
			12'd1222 : q <= 23'h362861; 
			12'd1223 : q <= 23'h242821; 
			12'd1224 : q <= 23'h34906d; 
			12'd1225 : q <= 23'h232481; 
			12'd1226 : q <= 23'h280846; 
			12'd1227 : q <= 23'h3048c1; 
			12'd1228 : q <= 23'h253c65; 
			12'd1229 : q <= 23'h349c25; 
			12'd1230 : q <= 23'h251043; 
			12'd1231 : q <= 23'h349028; 
			12'd1232 : q <= 23'h34986d; 
			12'd1233 : q <= 23'h230086; 
			12'd1234 : q <= 23'h380848; 
			12'd1235 : q <= 23'h338026; 
			12'd1236 : q <= 23'h380848; 
			12'd1237 : q <= 23'h2020c3; 
			12'd1238 : q <= 23'h263061; 
			12'd1239 : q <= 23'h34c422; 
			12'd1240 : q <= 23'h261821; 
			12'd1241 : q <= 23'h33a4c2; 
			12'd1242 : q <= 23'h261821; 
			12'd1243 : q <= 23'h339088; 
			12'd1244 : q <= 23'h36b0a1; 
			12'd1245 : q <= 23'h34ac41; 
			12'd1246 : q <= 23'h271c23; 
			12'd1247 : q <= 23'h329421; 
			12'd1248 : q <= 23'h369441; 
			12'd1249 : q <= 23'h329441; 
			12'd1250 : q <= 23'h34a441; 
			12'd1251 : q <= 23'h242841; 
			12'd1252 : q <= 23'h27c022; 
			12'd1253 : q <= 23'h21b441; 
			12'd1254 : q <= 23'h26bc21; 
			12'd1255 : q <= 23'h24b841; 
			12'd1256 : q <= 23'h3239c3; 
			12'd1257 : q <= 23'h33b881; 
			12'd1258 : q <= 23'h27c022; 
			12'd1259 : q <= 23'h224022; 
			12'd1260 : q <= 23'h38004d; 
			12'd1261 : q <= 23'h220426; 
			12'd1262 : q <= 23'h273863; 
			12'd1263 : q <= 23'h21b863; 
			12'd1264 : q <= 23'h274861; 
			12'd1265 : q <= 23'h21c861; 
			12'd1266 : q <= 23'h38004d; 
			12'd1267 : q <= 23'h31004d; 
			12'd1268 : q <= 23'h3530e2; 
			12'd1269 : q <= 23'h233c21; 
			12'd1270 : q <= 23'h252c83; 
			12'd1271 : q <= 23'h239821; 
			12'd1272 : q <= 23'h250903; 
			12'd1273 : q <= 23'h329461; 
			12'd1274 : q <= 23'h25b065; 
			12'd1275 : q <= 23'h233065; 
			12'd1276 : q <= 23'h359c22; 
			12'd1277 : q <= 23'h243481; 
			12'd1278 : q <= 23'h350821; 
			12'd1279 : q <= 23'h208849; 
			12'd1280 : q <= 23'h262886; 
			12'd1281 : q <= 23'h300822; 
			12'd1282 : q <= 23'h34b041; 
			12'd1283 : q <= 23'h342081; 
			12'd1284 : q <= 23'h359c22; 
			12'd1285 : q <= 23'h341c22; 
			12'd1286 : q <= 23'h359041; 
			12'd1287 : q <= 23'h249c23; 
			12'd1288 : q <= 23'h281c83; 
			12'd1289 : q <= 23'h201c83; 
			12'd1290 : q <= 23'h298825; 
			12'd1291 : q <= 23'h218864; 
			12'd1292 : q <= 23'h359041; 
			12'd1293 : q <= 23'h23bc21; 
			12'd1294 : q <= 23'h25c023; 
			12'd1295 : q <= 23'h244023; 
			12'd1296 : q <= 23'h270c21; 
			12'd1297 : q <= 23'h344041; 
			12'd1298 : q <= 23'h2644e2; 
			12'd1299 : q <= 23'h323d81; 
			12'd1300 : q <= 23'h358c22; 
			12'd1301 : q <= 23'h223441; 
			12'd1302 : q <= 23'h253883; 
			12'd1303 : q <= 23'h23b421; 
			12'd1304 : q <= 23'h25ace2; 
			12'd1305 : q <= 23'h33c8c2; 
			12'd1306 : q <= 23'h264821; 
			12'd1307 : q <= 23'h23c821; 
			12'd1308 : q <= 23'h264d01; 
			12'd1309 : q <= 23'h23bcc1; 
			12'd1310 : q <= 23'h253044; 
			12'd1311 : q <= 23'h322861; 
			12'd1312 : q <= 23'h34a842; 
			12'd1313 : q <= 23'h23804f; 
			12'd1314 : q <= 23'h36188e; 
			12'd1315 : q <= 23'h32c461; 
			12'd1316 : q <= 23'h360493; 
			12'd1317 : q <= 23'h218461; 
			12'd1318 : q <= 23'h253045; 
			12'd1319 : q <= 23'h243045; 
			12'd1320 : q <= 23'h262c21; 
			12'd1321 : q <= 23'h301062; 
			12'd1322 : q <= 23'h262c21; 
			12'd1323 : q <= 23'h23ac85; 
			12'd1324 : q <= 23'h262c21; 
			12'd1325 : q <= 23'h2138a1; 
			12'd1326 : q <= 23'h262c21; 
			12'd1327 : q <= 23'h23ac21; 
			12'd1328 : q <= 23'h373861; 
			12'd1329 : q <= 23'h31b861; 
			12'd1330 : q <= 23'h34bc41; 
			12'd1331 : q <= 23'h342061; 
			12'd1332 : q <= 23'h369861; 
			12'd1333 : q <= 23'h3028a1; 
			12'd1334 : q <= 23'h369861; 
			12'd1335 : q <= 23'h24b024; 
			12'd1336 : q <= 23'h261c21; 
			12'd1337 : q <= 23'h21c064; 
			12'd1338 : q <= 23'h351c41; 
			12'd1339 : q <= 23'h349c42; 
			12'd1340 : q <= 23'h263c84; 
			12'd1341 : q <= 23'h223886; 
			12'd1342 : q <= 23'h350022; 
			12'd1343 : q <= 23'h233c42; 
			12'd1344 : q <= 23'h369c2d; 
			12'd1345 : q <= 23'h331c2d; 
			12'd1346 : q <= 23'h34a463; 
			12'd1347 : q <= 23'h2228e6; 
			12'd1348 : q <= 23'h26b021; 
			12'd1349 : q <= 23'h233021; 
			12'd1350 : q <= 23'h252441; 
			12'd1351 : q <= 23'h219821; 
			12'd1352 : q <= 23'h281c61; 
			12'd1353 : q <= 23'h202662; 
			12'd1354 : q <= 23'h2508a1; 
			12'd1355 : q <= 23'h24a846; 
			12'd1356 : q <= 23'h264841; 
			12'd1357 : q <= 23'h209c62; 
			12'd1358 : q <= 23'h37004d; 
			12'd1359 : q <= 23'h32004d; 
			12'd1360 : q <= 23'h252504; 
			12'd1361 : q <= 23'h248c25; 
			12'd1362 : q <= 23'h359061; 
			12'd1363 : q <= 23'h331061; 
			12'd1364 : q <= 23'h3380ca; 
			12'd1365 : q <= 23'h33c8a1; 
			12'd1366 : q <= 23'h34ac41; 
			12'd1367 : q <= 23'h210c61; 
			12'd1368 : q <= 23'h243481; 
			12'd1369 : q <= 23'h233463; 
			12'd1370 : q <= 23'h259024; 
			12'd1371 : q <= 23'h241024; 
			12'd1372 : q <= 23'h249824; 
			12'd1373 : q <= 23'h333901; 
			12'd1374 : q <= 23'h353c24; 
			12'd1375 : q <= 23'h250831; 
			12'd1376 : q <= 23'h348041; 
			12'd1377 : q <= 23'h34bc24; 
			12'd1378 : q <= 23'h33b8e1; 
			12'd1379 : q <= 23'h34c023; 
			12'd1380 : q <= 23'h231d05; 
			12'd1381 : q <= 23'h212504; 
			12'd1382 : q <= 23'h274441; 
			12'd1383 : q <= 23'h224441; 
			12'd1384 : q <= 23'h253883; 
			12'd1385 : q <= 23'h233883; 
			12'd1386 : q <= 23'h353c21; 
			12'd1387 : q <= 23'h343c81; 
			12'd1388 : q <= 23'h260043; 
			12'd1389 : q <= 23'h201281; 
			12'd1390 : q <= 23'h280081; 
			12'd1391 : q <= 23'h214144; 
			12'd1392 : q <= 23'h291c25; 
			12'd1393 : q <= 23'h209c25; 
			12'd1394 : q <= 23'h37b062; 
			12'd1395 : q <= 23'h331042; 
			12'd1396 : q <= 23'h301e82; 
			12'd1397 : q <= 23'h200081; 
			12'd1398 : q <= 23'h3380c4; 
			12'd1399 : q <= 23'h20b8c1; 
			12'd1400 : q <= 23'h35a024; 
			12'd1401 : q <= 23'h340441; 
			12'd1402 : q <= 23'h343c81; 
			12'd1403 : q <= 23'h251922; 
			12'd1404 : q <= 23'h27b021; 
			12'd1405 : q <= 23'h231821; 
			12'd1406 : q <= 23'h369421; 
			12'd1407 : q <= 23'h214021; 
			12'd1408 : q <= 23'h361481; 
			12'd1409 : q <= 23'h3004e1; 
			12'd1410 : q <= 23'h24b062; 
			12'd1411 : q <= 23'h329441; 
			12'd1412 : q <= 23'h391441; 
			12'd1413 : q <= 23'h318902; 
			12'd1414 : q <= 23'h250943; 
			12'd1415 : q <= 23'h229c24; 
			12'd1416 : q <= 23'h3428a2; 
			12'd1417 : q <= 23'h2480cb; 
			12'd1418 : q <= 23'h268026; 
			12'd1419 : q <= 23'h20cc21; 
			12'd1420 : q <= 23'h292845; 
			12'd1421 : q <= 23'h322541; 
			12'd1422 : q <= 23'h373461; 
			12'd1423 : q <= 23'h202845; 
			12'd1424 : q <= 23'h391442; 
			12'd1425 : q <= 23'h331c21; 
			12'd1426 : q <= 23'h23a0e1; 
			12'd1427 : q <= 23'h301442; 
			12'd1428 : q <= 23'h360421; 
			12'd1429 : q <= 23'h230026; 
			12'd1430 : q <= 23'h3384ce; 
			12'd1431 : q <= 23'h241883; 
			12'd1432 : q <= 23'h24b062; 
			12'd1433 : q <= 23'h243062; 
			12'd1434 : q <= 23'h359c25; 
			12'd1435 : q <= 23'h341c25; 
			12'd1436 : q <= 23'h37002a; 
			12'd1437 : q <= 23'h223061; 
			12'd1438 : q <= 23'h390c26; 
			12'd1439 : q <= 23'h20b645; 
			12'd1440 : q <= 23'h37002a; 
			12'd1441 : q <= 23'h34bc41; 
			12'd1442 : q <= 23'h388c27; 
			12'd1443 : q <= 23'h32802a; 
			12'd1444 : q <= 23'h388c27; 
			12'd1445 : q <= 23'h202821; 
			12'd1446 : q <= 23'h29042a; 
			12'd1447 : q <= 23'h20842a; 
			12'd1448 : q <= 23'h35c024; 
			12'd1449 : q <= 23'h31a023; 
			12'd1450 : q <= 23'h260023; 
			12'd1451 : q <= 23'h238023; 
			12'd1452 : q <= 23'h388c27; 
			12'd1453 : q <= 23'h310c27; 
			12'd1454 : q <= 23'h380450; 
			12'd1455 : q <= 23'h310450; 
			12'd1456 : q <= 23'h250104; 
			12'd1457 : q <= 23'h3324a1; 
			12'd1458 : q <= 23'h351c23; 
			12'd1459 : q <= 23'h342481; 
			12'd1460 : q <= 23'h249824; 
			12'd1461 : q <= 23'h329ca1; 
			12'd1462 : q <= 23'h3414e3; 
			12'd1463 : q <= 23'h209d02; 
			12'd1464 : q <= 23'h233501; 
			12'd1465 : q <= 23'h343061; 
			12'd1466 : q <= 23'h2594e5; 
			12'd1467 : q <= 23'h223461; 
			12'd1468 : q <= 23'h35ac41; 
			12'd1469 : q <= 23'h322ce2; 
			12'd1470 : q <= 23'h33acc1; 
			12'd1471 : q <= 23'h24b041; 
			12'd1472 : q <= 23'h301e82; 
			12'd1473 : q <= 23'h341041; 
			12'd1474 : q <= 23'h35ac41; 
			12'd1475 : q <= 23'h33ac41; 
			12'd1476 : q <= 23'h35c024; 
			12'd1477 : q <= 23'h349c23; 
			12'd1478 : q <= 23'h214204; 
			12'd1479 : q <= 23'h2041e1; 
			12'd1480 : q <= 23'h3798a2; 
			12'd1481 : q <= 23'h251424; 
			12'd1482 : q <= 23'h343122; 
			12'd1483 : q <= 23'h33cca1; 
			12'd1484 : q <= 23'h35c024; 
			12'd1485 : q <= 23'h204682; 
			12'd1486 : q <= 23'h35c024; 
			12'd1487 : q <= 23'h344024; 
			12'd1488 : q <= 23'h34c461; 
			12'd1489 : q <= 23'h243883; 
			12'd1490 : q <= 23'h34a844; 
			12'd1491 : q <= 23'h344881; 
			12'd1492 : q <= 23'h26c881; 
			12'd1493 : q <= 23'h20cd01; 
			12'd1494 : q <= 23'h37944f; 
			12'd1495 : q <= 23'h24a441; 
			12'd1496 : q <= 23'h249423; 
			12'd1497 : q <= 23'h31944f; 
			12'd1498 : q <= 23'h2584e4; 
			12'd1499 : q <= 23'h211048; 
			12'd1500 : q <= 23'h262866; 
			12'd1501 : q <= 23'h2214a6; 
			12'd1502 : q <= 23'h34bc41; 
			12'd1503 : q <= 23'h329441; 
			12'd1504 : q <= 23'h270845; 
			12'd1505 : q <= 23'h3314e1; 
			12'd1506 : q <= 23'h258121; 
			12'd1507 : q <= 23'h200121; 
			12'd1508 : q <= 23'h27b443; 
			12'd1509 : q <= 23'h21b443; 
			12'd1510 : q <= 23'h253c43; 
			12'd1511 : q <= 23'h22a4a5; 
			12'd1512 : q <= 23'h269041; 
			12'd1513 : q <= 23'h253068; 
			12'd1514 : q <= 23'h270845; 
			12'd1515 : q <= 23'h24ac21; 
			12'd1516 : q <= 23'h352424; 
			12'd1517 : q <= 23'h21ac69; 
			12'd1518 : q <= 23'h270845; 
			12'd1519 : q <= 23'h220845; 
			12'd1520 : q <= 23'h269041; 
			12'd1521 : q <= 23'h303cc1; 
			12'd1522 : q <= 23'h269041; 
			12'd1523 : q <= 23'h338422; 
			12'd1524 : q <= 23'h269041; 
			12'd1525 : q <= 23'h229041; 
			12'd1526 : q <= 23'h270026; 
			12'd1527 : q <= 23'h33802a; 
			12'd1528 : q <= 23'h219224; 
			12'd1529 : q <= 23'h201a82; 
			12'd1530 : q <= 23'h220c82; 
			12'd1531 : q <= 23'h343081; 
			12'd1532 : q <= 23'h229c62; 
			12'd1533 : q <= 23'h341883; 
			12'd1534 : q <= 23'h244422; 
			12'd1535 : q <= 23'h341487; 
			12'd1536 : q <= 23'h220845; 
			12'd1537 : q <= 23'h218621; 
			12'd1538 : q <= 23'h311e05; 
			12'd1539 : q <= 23'h278ca1; 
			12'd1540 : q <= 23'h250c22; 
			12'd1541 : q <= 23'h322a05; 
			12'd1542 : q <= 23'h23c0a3; 
			12'd1543 : q <= 23'h359c22; 
			12'd1544 : q <= 23'h348c21; 
			12'd1545 : q <= 23'h34c461; 
			12'd1546 : q <= 23'h200ca1; 
			12'd1547 : q <= 23'h361881; 
			12'd1548 : q <= 23'h329c81; 
			12'd1549 : q <= 23'h23b0c7; 
			12'd1550 : q <= 23'h200085; 
			12'd1551 : q <= 23'h350422; 
			12'd1552 : q <= 23'h348422; 
			12'd1553 : q <= 23'h361461; 
			12'd1554 : q <= 23'h23b0c8; 
			12'd1555 : q <= 23'h361461; 
			12'd1556 : q <= 23'h311442; 
			12'd1557 : q <= 23'h3714c3; 
			12'd1558 : q <= 23'h329461; 
			12'd1559 : q <= 23'h354422; 
			12'd1560 : q <= 23'h329841; 
			12'd1561 : q <= 23'h36b462; 
			12'd1562 : q <= 23'h21c443; 
			12'd1563 : q <= 23'h2710c1; 
			12'd1564 : q <= 23'h202601; 
			12'd1565 : q <= 23'h2710c1; 
			12'd1566 : q <= 23'h3008a2; 
			12'd1567 : q <= 23'h361881; 
			12'd1568 : q <= 23'h323462; 
			12'd1569 : q <= 23'h361881; 
			12'd1570 : q <= 23'h349821; 
			12'd1571 : q <= 23'h361881; 
			12'd1572 : q <= 23'h233106; 
			12'd1573 : q <= 23'h361881; 
			12'd1574 : q <= 23'h343062; 
			12'd1575 : q <= 23'h361881; 
			12'd1576 : q <= 23'h321881; 
			12'd1577 : q <= 23'h349862; 
			12'd1578 : q <= 23'h323021; 
			12'd1579 : q <= 23'h273066; 
			12'd1580 : q <= 23'h340027; 
			12'd1581 : q <= 23'h352023; 
			12'd1582 : q <= 23'h34a023; 
			12'd1583 : q <= 23'h32ad61; 
			12'd1584 : q <= 23'h251ca1; 
			12'd1585 : q <= 23'h351c22; 
			12'd1586 : q <= 23'h349c22; 
			12'd1587 : q <= 23'h25a442; 
			12'd1588 : q <= 23'h23a442; 
			12'd1589 : q <= 23'h273042; 
			12'd1590 : q <= 23'h341c22; 
			12'd1591 : q <= 23'h3748c1; 
			12'd1592 : q <= 23'h2214c6; 
			12'd1593 : q <= 23'h252484; 
			12'd1594 : q <= 23'h3290a4; 
			12'd1595 : q <= 23'h268841; 
			12'd1596 : q <= 23'h223441; 
			12'd1597 : q <= 23'h343881; 
			12'd1598 : q <= 23'h34b841; 
			12'd1599 : q <= 23'h36b041; 
			12'd1600 : q <= 23'h23b042; 
			12'd1601 : q <= 23'h25ac21; 
			12'd1602 : q <= 23'h34c422; 
			12'd1603 : q <= 23'h25ac21; 
			12'd1604 : q <= 23'h3048c1; 
			12'd1605 : q <= 23'h25ac21; 
			12'd1606 : q <= 23'h242c21; 
			12'd1607 : q <= 23'h261484; 
			12'd1608 : q <= 23'h221484; 
			12'd1609 : q <= 23'h268841; 
			12'd1610 : q <= 23'h228841; 
			12'd1611 : q <= 23'h260041; 
			12'd1612 : q <= 23'h343021; 
			12'd1613 : q <= 23'h252c44; 
			12'd1614 : q <= 23'h24a841; 
			12'd1615 : q <= 23'h21cde1; 
			12'd1616 : q <= 23'h211826; 
			12'd1617 : q <= 23'h34a441; 
			12'd1618 : q <= 23'h342822; 
			12'd1619 : q <= 23'h362c21; 
			12'd1620 : q <= 23'h33ac21; 
			12'd1621 : q <= 23'h258841; 
			12'd1622 : q <= 23'h323441; 
			12'd1623 : q <= 23'h3404c3; 
			12'd1624 : q <= 23'h23844e; 
			12'd1625 : q <= 23'h2440c3; 
			12'd1626 : q <= 23'h33c4c3; 
			12'd1627 : q <= 23'h24c443; 
			12'd1628 : q <= 23'h24c024; 
			12'd1629 : q <= 23'h34bc41; 
			12'd1630 : q <= 23'h34a844; 
			12'd1631 : q <= 23'h362861; 
			12'd1632 : q <= 23'h210448; 
			12'd1633 : q <= 23'h260461; 
			12'd1634 : q <= 23'h20a987; 
			12'd1635 : q <= 23'h253041; 
			12'd1636 : q <= 23'h20a4a1; 
			12'd1637 : q <= 23'h344081; 
			12'd1638 : q <= 23'h332501; 
			12'd1639 : q <= 23'h34c0a1; 
			12'd1640 : q <= 23'h342081; 
			12'd1641 : q <= 23'h23a0c1; 
			12'd1642 : q <= 23'h229c81; 
			12'd1643 : q <= 23'h362861; 
			12'd1644 : q <= 23'h222081; 
			12'd1645 : q <= 23'h3714c3; 
			12'd1646 : q <= 23'h32a423; 
			12'd1647 : q <= 23'h362861; 
			12'd1648 : q <= 23'h3014c3; 
			12'd1649 : q <= 23'h390c26; 
			12'd1650 : q <= 23'h308c26; 
			12'd1651 : q <= 23'h28bc21; 
			12'd1652 : q <= 23'h232443; 
			12'd1653 : q <= 23'h362861; 
			12'd1654 : q <= 23'h32a861; 
			12'd1655 : q <= 23'h261464; 
			12'd1656 : q <= 23'h229464; 
			12'd1657 : q <= 23'h281083; 
			12'd1658 : q <= 23'h318054; 
			12'd1659 : q <= 23'h36ac22; 
			12'd1660 : q <= 23'h332c22; 
			12'd1661 : q <= 23'h359041; 
			12'd1662 : q <= 23'h220083; 
			12'd1663 : q <= 23'h278025; 
			12'd1664 : q <= 23'h328422; 
			12'd1665 : q <= 23'h34804f; 
			12'd1666 : q <= 23'h33ac21; 
			12'd1667 : q <= 23'h368024; 
			12'd1668 : q <= 23'h339041; 
			12'd1669 : q <= 23'h262061; 
			12'd1670 : q <= 23'h201083; 
			12'd1671 : q <= 23'h262061; 
			12'd1672 : q <= 23'h314461; 
			12'd1673 : q <= 23'h282065; 
			12'd1674 : q <= 23'h2028a1; 
			12'd1675 : q <= 23'h26ac21; 
			12'd1676 : q <= 23'h31c061; 
			12'd1677 : q <= 23'h262061; 
			12'd1678 : q <= 23'h22a061; 
			12'd1679 : q <= 23'h34a123; 
			12'd1680 : q <= 23'h330027; 
			12'd1681 : q <= 23'h348885; 
			12'd1682 : q <= 23'h232c21; 
			12'd1683 : q <= 23'h27c061; 
			12'd1684 : q <= 23'h214061; 
			12'd1685 : q <= 23'h28b064; 
			12'd1686 : q <= 23'h33a0a6; 
			12'd1687 : q <= 23'h3408d1; 
			12'd1688 : q <= 23'h238441; 
			12'd1689 : q <= 23'h348885; 
			12'd1690 : q <= 23'h338885; 
			12'd1691 : q <= 23'h2524c2; 
			12'd1692 : q <= 23'h22bc61; 
			12'd1693 : q <= 23'h353c41; 
			12'd1694 : q <= 23'h203541; 
			12'd1695 : q <= 23'h2524c4; 
			12'd1696 : q <= 23'h244063; 
			12'd1697 : q <= 23'h253441; 
			12'd1698 : q <= 23'h24b021; 
			12'd1699 : q <= 23'h25ace2; 
			12'd1700 : q <= 23'h241881; 
			12'd1701 : q <= 23'h362843; 
			12'd1702 : q <= 23'h213c21; 
			12'd1703 : q <= 23'h282066; 
			12'd1704 : q <= 23'h20a066; 
			12'd1705 : q <= 23'h36004a; 
			12'd1706 : q <= 23'h22ac82; 
			12'd1707 : q <= 23'h274082; 
			12'd1708 : q <= 23'h349c46; 
			12'd1709 : q <= 23'h25084a; 
			12'd1710 : q <= 23'h240449; 
			12'd1711 : q <= 23'h264c21; 
			12'd1712 : q <= 23'h218849; 
			12'd1713 : q <= 23'h349444; 
			12'd1714 : q <= 23'h249842; 
			12'd1715 : q <= 23'h272444; 
			12'd1716 : q <= 23'h23b0a6; 
			12'd1717 : q <= 23'h272443; 
			12'd1718 : q <= 23'h222443; 
			12'd1719 : q <= 23'h26bca2; 
			12'd1720 : q <= 23'h23c822; 
			12'd1721 : q <= 23'h2590c1; 
			12'd1722 : q <= 23'h310a02; 
			12'd1723 : q <= 23'h2590c1; 
			12'd1724 : q <= 23'h323141; 
			12'd1725 : q <= 23'h2590c1; 
			12'd1726 : q <= 23'h2190c1; 
			12'd1727 : q <= 23'h280047; 
			12'd1728 : q <= 23'h304122; 
			12'd1729 : q <= 23'h34c461; 
			12'd1730 : q <= 23'h331842; 
			12'd1731 : q <= 23'h37b021; 
			12'd1732 : q <= 23'h329841; 
			12'd1733 : q <= 23'h252841; 
			12'd1734 : q <= 23'h228443; 
			12'd1735 : q <= 23'h280047; 
			12'd1736 : q <= 23'h250141; 
			12'd1737 : q <= 23'h37b021; 
			12'd1738 : q <= 23'h309024; 
			12'd1739 : q <= 23'h381462; 
			12'd1740 : q <= 23'h309462; 
			12'd1741 : q <= 23'h2608c3; 
			12'd1742 : q <= 23'h342c81; 
			12'd1743 : q <= 23'h2588e3; 
			12'd1744 : q <= 23'h34b041; 
			12'd1745 : q <= 23'h37b841; 
			12'd1746 : q <= 23'h343481; 
			12'd1747 : q <= 23'h37b021; 
			12'd1748 : q <= 23'h23b8a1; 
			12'd1749 : q <= 23'h33b4c1; 
			12'd1750 : q <= 23'h22b482; 
			12'd1751 : q <= 23'h361023; 
			12'd1752 : q <= 23'h339023; 
			12'd1753 : q <= 23'h389426; 
			12'd1754 : q <= 23'h339887; 
			12'd1755 : q <= 23'h389426; 
			12'd1756 : q <= 23'h31b841; 
			12'd1757 : q <= 23'h389426; 
			12'd1758 : q <= 23'h311426; 
			12'd1759 : q <= 23'h33a4c1; 
			12'd1760 : q <= 23'h222487; 
			12'd1761 : q <= 23'h263101; 
			12'd1762 : q <= 23'h203101; 
			12'd1763 : q <= 23'h34b841; 
			12'd1764 : q <= 23'h2228c2; 
			12'd1765 : q <= 23'h350c27; 
			12'd1766 : q <= 23'h340825; 
			12'd1767 : q <= 23'h25b043; 
			12'd1768 : q <= 23'h349c26; 
			12'd1769 : q <= 23'h279481; 
			12'd1770 : q <= 23'h349c23; 
			12'd1771 : q <= 23'h2710c2; 
			12'd1772 : q <= 23'h34c041; 
			12'd1773 : q <= 23'h37b841; 
			12'd1774 : q <= 23'h349c2a; 
			12'd1775 : q <= 23'h35b042; 
			12'd1776 : q <= 23'h242841; 
			12'd1777 : q <= 23'h252841; 
			12'd1778 : q <= 23'h242841; 
			12'd1779 : q <= 23'h269c21; 
			12'd1780 : q <= 23'h229c21; 
			12'd1781 : q <= 23'h37002e; 
			12'd1782 : q <= 23'h32802e; 
			12'd1783 : q <= 23'h37102e; 
			12'd1784 : q <= 23'h34bc41; 
			12'd1785 : q <= 23'h343c81; 
			12'd1786 : q <= 23'h328830; 
			12'd1787 : q <= 23'h239d05; 
			12'd1788 : q <= 23'h333ce1; 
			12'd1789 : q <= 23'h2708a6; 
			12'd1790 : q <= 23'h232101; 
			12'd1791 : q <= 23'h244083; 
			12'd1792 : q <= 23'h331c21; 
			12'd1793 : q <= 23'h381082; 
			12'd1794 : q <= 23'h231841; 
			12'd1795 : q <= 23'h381082; 
			12'd1796 : q <= 23'h301082; 
			12'd1797 : q <= 23'h249826; 
			12'd1798 : q <= 23'h21a4c5; 
			12'd1799 : q <= 23'h249426; 
			12'd1800 : q <= 23'h31b841; 
			12'd1801 : q <= 23'h26b861; 
			12'd1802 : q <= 23'h2140a2; 
			12'd1803 : q <= 23'h2518a3; 
			12'd1804 : q <= 23'h33bc21; 
			12'd1805 : q <= 23'h3744c1; 
			12'd1806 : q <= 23'h329461; 
			12'd1807 : q <= 23'h339541; 
			12'd1808 : q <= 23'h2018a2; 
			12'd1809 : q <= 23'h36b863; 
			12'd1810 : q <= 23'h323863; 
			12'd1811 : q <= 23'h249c21; 
			12'd1812 : q <= 23'h338051; 
			12'd1813 : q <= 23'h250c63; 
			12'd1814 : q <= 23'h3388a4; 
			12'd1815 : q <= 23'h260881; 
			12'd1816 : q <= 23'h340c62; 
			12'd1817 : q <= 23'h24c841; 
			12'd1818 : q <= 23'h20802e; 
			12'd1819 : q <= 23'h3604e1; 
			12'd1820 : q <= 23'h20bc21; 
			12'd1821 : q <= 23'h27b024; 
			12'd1822 : q <= 23'h3084e1; 
			12'd1823 : q <= 23'h27b024; 
			12'd1824 : q <= 23'h230086; 
			12'd1825 : q <= 23'h331103; 
			12'd1826 : q <= 23'h228c41; 
			12'd1827 : q <= 23'h283863; 
			12'd1828 : q <= 23'h204541; 
			12'd1829 : q <= 23'h258c23; 
			12'd1830 : q <= 23'h243062; 
			12'd1831 : q <= 23'h251c6d; 
			12'd1832 : q <= 23'h253ca5; 
			12'd1833 : q <= 23'h25104a; 
			12'd1834 : q <= 23'h231c21; 
			12'd1835 : q <= 23'h250c67; 
			12'd1836 : q <= 23'h238c67; 
			12'd1837 : q <= 23'h339cc5; 
			12'd1838 : q <= 23'h22c443; 
			12'd1839 : q <= 23'h2738c3; 
			12'd1840 : q <= 23'h203542; 
			12'd1841 : q <= 23'h2594e1; 
			12'd1842 : q <= 23'h2088a6; 
			12'd1843 : q <= 23'h3309c1; 
			12'd1844 : q <= 23'h344441; 
			12'd1845 : q <= 23'h354422; 
			12'd1846 : q <= 23'h22bc41; 
			12'd1847 : q <= 23'h354021; 
			12'd1848 : q <= 23'h244042; 
			12'd1849 : q <= 23'h233903; 
			12'd1850 : q <= 23'h2138a1; 
			12'd1851 : q <= 23'h283863; 
			12'd1852 : q <= 23'h33a4c4; 
			12'd1853 : q <= 23'h283863; 
			12'd1854 : q <= 23'h301022; 
			12'd1855 : q <= 23'h22a9ea; 
			12'd1856 : q <= 23'h20b863; 
			12'd1857 : q <= 23'h253843; 
			12'd1858 : q <= 23'h242c21; 
			12'd1859 : q <= 23'h354422; 
			12'd1860 : q <= 23'h34c422; 
			12'd1861 : q <= 23'h273843; 
			12'd1862 : q <= 23'h223843; 
			12'd1863 : q <= 23'h273823; 
			12'd1864 : q <= 23'h22b823; 
			12'd1865 : q <= 23'h3390c4; 
			12'd1866 : q <= 23'h321c82; 
			12'd1867 : q <= 23'h358c2d; 
			12'd1868 : q <= 23'h340c2d; 
			12'd1869 : q <= 23'h3524c1; 
			12'd1870 : q <= 23'h322c22; 
			12'd1871 : q <= 23'h283064; 
			12'd1872 : q <= 23'h349845; 
			12'd1873 : q <= 23'h28ac27; 
			12'd1874 : q <= 23'h23b482; 
			12'd1875 : q <= 23'h332901; 
			12'd1876 : q <= 23'h321081; 
			12'd1877 : q <= 23'h359081; 
			12'd1878 : q <= 23'h30a224; 
			12'd1879 : q <= 23'h359081; 
			12'd1880 : q <= 23'h3224c1; 
			12'd1881 : q <= 23'h3610a1; 
			12'd1882 : q <= 23'h212c27; 
			12'd1883 : q <= 23'h283024; 
			12'd1884 : q <= 23'h322561; 
			12'd1885 : q <= 23'h263461; 
			12'd1886 : q <= 23'h333881; 
			12'd1887 : q <= 23'h353023; 
			12'd1888 : q <= 23'h329061; 
			12'd1889 : q <= 23'h349441; 
			12'd1890 : q <= 23'h300e01; 
			12'd1891 : q <= 23'h283024; 
			12'd1892 : q <= 23'h21b024; 
			12'd1893 : q <= 23'h373c62; 
			12'd1894 : q <= 23'h31bc62; 
			12'd1895 : q <= 23'h2594a1; 
			12'd1896 : q <= 23'h2145c3; 
			12'd1897 : q <= 23'h353c21; 
			12'd1898 : q <= 23'h224021; 
			12'd1899 : q <= 23'h351c41; 
			12'd1900 : q <= 23'h204541; 
			12'd1901 : q <= 23'h369c21; 
			12'd1902 : q <= 23'h34b422; 
			12'd1903 : q <= 23'h368823; 
			12'd1904 : q <= 23'h21c821; 
			12'd1905 : q <= 23'h354024; 
			12'd1906 : q <= 23'h331c21; 
			12'd1907 : q <= 23'h2688a1; 
			12'd1908 : q <= 23'h23b861; 
			12'd1909 : q <= 23'h360c24; 
			12'd1910 : q <= 23'h32b486; 
			12'd1911 : q <= 23'h2730a1; 
			12'd1912 : q <= 23'h213ce2; 
			12'd1913 : q <= 23'h251ce1; 
			12'd1914 : q <= 23'h20b081; 
			12'd1915 : q <= 23'h38004e; 
			12'd1916 : q <= 23'h323021; 
			12'd1917 : q <= 23'h38004e; 
			12'd1918 : q <= 23'h312827; 
			12'd1919 : q <= 23'h243521; 
			12'd1920 : q <= 23'h251941; 
			12'd1921 : q <= 23'h241044; 
			12'd1922 : q <= 23'h200441; 
			12'd1923 : q <= 23'h329943; 
			12'd1924 : q <= 23'h27884a; 
			12'd1925 : q <= 23'h248827; 
			12'd1926 : q <= 23'h359081; 
			12'd1927 : q <= 23'h331061; 
			12'd1928 : q <= 23'h27b022; 
			12'd1929 : q <= 23'h23a864; 
			12'd1930 : q <= 23'h27b023; 
			12'd1931 : q <= 23'h33c8c1; 
			12'd1932 : q <= 23'h278c28; 
			12'd1933 : q <= 23'h223023; 
			12'd1934 : q <= 23'h2608a1; 
			12'd1935 : q <= 23'h234841; 
			12'd1936 : q <= 23'h251105; 
			12'd1937 : q <= 23'h232825; 
			12'd1938 : q <= 23'h34a0a2; 
			12'd1939 : q <= 23'h3320a2; 
			12'd1940 : q <= 23'h349c62; 
			12'd1941 : q <= 23'h249c82; 
			12'd1942 : q <= 23'h34b041; 
			12'd1943 : q <= 23'h308601; 
			12'd1944 : q <= 23'h258ce1; 
			12'd1945 : q <= 23'h329d46; 
			12'd1946 : q <= 23'h391022; 
			12'd1947 : q <= 23'h343821; 
			12'd1948 : q <= 23'h31c1c2; 
			12'd1949 : q <= 23'h308824; 
			12'd1950 : q <= 23'h2608a1; 
			12'd1951 : q <= 23'h2188a1; 
			12'd1952 : q <= 23'h353841; 
			12'd1953 : q <= 23'h343841; 
			12'd1954 : q <= 23'h373441; 
			12'd1955 : q <= 23'h338c41; 
			12'd1956 : q <= 23'h2518a2; 
			12'd1957 : q <= 23'h24c023; 
			12'd1958 : q <= 23'h25b021; 
			12'd1959 : q <= 23'h323441; 
			12'd1960 : q <= 23'h3718c2; 
			12'd1961 : q <= 23'h344841; 
			12'd1962 : q <= 23'h381882; 
			12'd1963 : q <= 23'h301882; 
			12'd1964 : q <= 23'h271823; 
			12'd1965 : q <= 23'h242481; 
			12'd1966 : q <= 23'h343481; 
			12'd1967 : q <= 23'h32b942; 
			12'd1968 : q <= 23'h25b421; 
			12'd1969 : q <= 23'h244081; 
			12'd1970 : q <= 23'h252484; 
			12'd1971 : q <= 23'h23b043; 
			12'd1972 : q <= 23'h35ac21; 
			12'd1973 : q <= 23'h249c25; 
			12'd1974 : q <= 23'h350046; 
			12'd1975 : q <= 23'h31b442; 
			12'd1976 : q <= 23'h283421; 
			12'd1977 : q <= 23'h20b863; 
			12'd1978 : q <= 23'h370426; 
			12'd1979 : q <= 23'h242441; 
			12'd1980 : q <= 23'h352423; 
			12'd1981 : q <= 23'h342061; 
			12'd1982 : q <= 23'h270023; 
			12'd1983 : q <= 23'h3380c9; 
			12'd1984 : q <= 23'h25944f; 
			12'd1985 : q <= 23'h23944f; 
			12'd1986 : q <= 23'h270023; 
			12'd1987 : q <= 23'h228023; 
			12'd1988 : q <= 23'h263021; 
			12'd1989 : q <= 23'h23b021; 
			12'd1990 : q <= 23'h368024; 
			12'd1991 : q <= 23'h323061; 
			12'd1992 : q <= 23'h262081; 
			12'd1993 : q <= 23'h34a822; 
			12'd1994 : q <= 23'h352422; 
			12'd1995 : q <= 23'h34a422; 
			12'd1996 : q <= 23'h368024; 
			12'd1997 : q <= 23'h330024; 
			12'd1998 : q <= 23'h2538c2; 
			12'd1999 : q <= 23'h343841; 
			12'd2000 : q <= 23'h253864; 
			12'd2001 : q <= 23'h242844; 
			12'd2002 : q <= 23'h35a021; 
			12'd2003 : q <= 23'h24bc23; 
			12'd2004 : q <= 23'h35a021; 
			12'd2005 : q <= 23'h342021; 
			12'd2006 : q <= 23'h22a5e7; 
			12'd2007 : q <= 23'h210425; 
			12'd2008 : q <= 23'h373c41; 
			12'd2009 : q <= 23'h319c23; 
			12'd2010 : q <= 23'h389461; 
			12'd2011 : q <= 23'h301461; 
			12'd2012 : q <= 23'h281461; 
			12'd2013 : q <= 23'h344c81; 
			12'd2014 : q <= 23'h263842; 
			12'd2015 : q <= 23'h31c021; 
			12'd2016 : q <= 23'h25c064; 
			12'd2017 : q <= 23'h31a82a; 
			12'd2018 : q <= 23'h262024; 
			12'd2019 : q <= 23'h23a024; 
			12'd2020 : q <= 23'h253823; 
			12'd2021 : q <= 23'h2504a3; 
			12'd2022 : q <= 23'h359c22; 
			12'd2023 : q <= 23'h341862; 
			12'd2024 : q <= 23'h24a441; 
			12'd2025 : q <= 23'h212d03; 
			12'd2026 : q <= 23'h269c21; 
			12'd2027 : q <= 23'h349841; 
			12'd2028 : q <= 23'h351c22; 
			12'd2029 : q <= 23'h229d06; 
			12'd2030 : q <= 23'h269841; 
			12'd2031 : q <= 23'h229841; 
			12'd2032 : q <= 23'h361461; 
			12'd2033 : q <= 23'h323c41; 
			12'd2034 : q <= 23'h361461; 
			12'd2035 : q <= 23'h329461; 
			12'd2036 : q <= 23'h253823; 
			12'd2037 : q <= 23'h34b822; 
			12'd2038 : q <= 23'h359446; 
			12'd2039 : q <= 23'h339446; 
			12'd2040 : q <= 23'h26b821; 
			12'd2041 : q <= 23'h200d41; 
			12'd2042 : q <= 23'h26b821; 
			12'd2043 : q <= 23'h229c21; 
			12'd2044 : q <= 23'h269427; 
			12'd2045 : q <= 23'h233821; 
			12'd2046 : q <= 23'h360027; 
			12'd2047 : q <= 23'h200c28; 
			12'd2048 : q <= 23'h360027; 
			12'd2049 : q <= 23'h338027; 
			12'd2050 : q <= 23'h25c084; 
			12'd2051 : q <= 23'h22c084; 
			12'd2052 : q <= 23'h269427; 
			12'd2053 : q <= 23'h231427; 
			12'd2054 : q <= 23'h293447; 
			12'd2055 : q <= 23'h233062; 
			12'd2056 : q <= 23'h272021; 
			12'd2057 : q <= 23'h200523; 
			12'd2058 : q <= 23'h272021; 
			12'd2059 : q <= 23'h203447; 
			12'd2060 : q <= 23'h39002c; 
			12'd2061 : q <= 23'h301e41; 
			12'd2062 : q <= 23'h2321c8; 
			12'd2063 : q <= 23'h30802c; 
			12'd2064 : q <= 23'h370027; 
			12'd2065 : q <= 23'h22a021; 
			12'd2066 : q <= 23'h3718c2; 
			12'd2067 : q <= 23'h22a0e1; 
			12'd2068 : q <= 23'h3424c3; 
			12'd2069 : q <= 23'h339041; 
			12'd2070 : q <= 23'h280062; 
			12'd2071 : q <= 23'h309a44; 
			12'd2072 : q <= 23'h319a24; 
			12'd2073 : q <= 23'h32bce1; 
			12'd2074 : q <= 23'h353c21; 
			12'd2075 : q <= 23'h31bc61; 
			12'd2076 : q <= 23'h3718c2; 
			12'd2077 : q <= 23'h3018c2; 
			12'd2078 : q <= 23'h361881; 
			12'd2079 : q <= 23'h321881; 
			12'd2080 : q <= 23'h390842; 
			12'd2081 : q <= 23'h250449; 
			12'd2082 : q <= 23'h231882; 
			12'd2083 : q <= 23'h231441; 
			12'd2084 : q <= 23'h351841; 
			12'd2085 : q <= 23'h349821; 
			12'd2086 : q <= 23'h24ac41; 
			12'd2087 : q <= 23'h302481; 
			12'd2088 : q <= 23'h230d03; 
			12'd2089 : q <= 23'h208062; 
			12'd2090 : q <= 23'h370027; 
			12'd2091 : q <= 23'h24c441; 
			12'd2092 : q <= 23'h25a4c5; 
			12'd2093 : q <= 23'h202e61; 
			12'd2094 : q <= 23'h34a103; 
			12'd2095 : q <= 23'h328027; 
			12'd2096 : q <= 23'h251846; 
			12'd2097 : q <= 23'h2010c2; 
			12'd2098 : q <= 23'h344081; 
			12'd2099 : q <= 23'h348027; 
			12'd2100 : q <= 23'h351424; 
			12'd2101 : q <= 23'h349424; 
			12'd2102 : q <= 23'h349841; 
			12'd2103 : q <= 23'h23b842; 
			12'd2104 : q <= 23'h27b843; 
			12'd2105 : q <= 23'h23b024; 
			12'd2106 : q <= 23'h288024; 
			12'd2107 : q <= 23'h210024; 
			12'd2108 : q <= 23'h3309c1; 
			12'd2109 : q <= 23'h23b865; 
			12'd2110 : q <= 23'h24bc41; 
			12'd2111 : q <= 23'h23acc4; 
			12'd2112 : q <= 23'h24a863; 
			12'd2113 : q <= 23'h33b861; 
			12'd2114 : q <= 23'h24a841; 
			12'd2115 : q <= 23'h3304c2; 
			12'd2116 : q <= 23'h23a0c7; 
			12'd2117 : q <= 23'h33a4c1; 
			12'd2118 : q <= 23'h249c22; 
			12'd2119 : q <= 23'h250c29; 
			12'd2120 : q <= 23'h393c41; 
			12'd2121 : q <= 23'h342c21; 
			12'd2122 : q <= 23'h35a024; 
			12'd2123 : q <= 23'h343826; 
			12'd2124 : q <= 23'h35a024; 
			12'd2125 : q <= 23'h342024; 
			12'd2126 : q <= 23'h33b0c3; 
			12'd2127 : q <= 23'h303c41; 
			12'd2128 : q <= 23'h25b421; 
			12'd2129 : q <= 23'h240c83; 
			12'd2130 : q <= 23'h201146; 
			12'd2131 : q <= 23'h34bc21; 
			12'd2132 : q <= 23'h343c81; 
			12'd2133 : q <= 23'h2045c2; 
			12'd2134 : q <= 23'h20c643; 
			12'd2135 : q <= 23'h2000a3;
			default	 : q <= 23'h000000;
		endcase	
	end
	assign out = q;
endmodule